VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_96x4096_1rw
  FOREIGN sram_96x4096_1rw 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 747.080 BY 572.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.185 0.070 3.255 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.825 0.070 6.895 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.105 0.070 14.175 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.745 0.070 17.815 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.025 0.070 25.095 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.665 0.070 28.735 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.945 0.070 36.015 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.405 0.070 41.475 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.505 0.070 50.575 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.785 0.070 57.855 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.425 0.070 61.495 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.245 0.070 63.315 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.705 0.070 68.775 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.345 0.070 72.415 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.625 0.070 79.695 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.265 0.070 83.335 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.085 0.070 85.155 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.725 0.070 88.795 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.545 0.070 90.615 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.185 0.070 94.255 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.005 0.070 96.075 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.825 0.070 97.895 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.465 0.070 101.535 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.105 0.070 105.175 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.925 0.070 106.995 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.565 0.070 110.635 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.385 0.070 112.455 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.205 0.070 114.275 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.025 0.070 116.095 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.845 0.070 117.915 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.665 0.070 119.735 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.305 0.070 123.375 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.125 0.070 125.195 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.945 0.070 127.015 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.585 0.070 130.655 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.405 0.070 132.475 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.225 0.070 134.295 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.045 0.070 136.115 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.865 0.070 137.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.685 0.070 139.755 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.505 0.070 141.575 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.145 0.070 145.215 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.965 0.070 147.035 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.785 0.070 148.855 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.425 0.070 152.495 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.065 0.070 156.135 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.885 0.070 157.955 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.705 0.070 159.775 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.525 0.070 161.595 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.345 0.070 163.415 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.985 0.070 167.055 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.805 0.070 168.875 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.625 0.070 170.695 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.445 0.070 172.515 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.265 0.070 174.335 ;
    END
  END w_mask_in[95]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.745 0.070 178.815 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.565 0.070 180.635 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.385 0.070 182.455 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.205 0.070 184.275 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.025 0.070 186.095 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.845 0.070 187.915 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.665 0.070 189.735 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.485 0.070 191.555 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.305 0.070 193.375 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.125 0.070 195.195 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.945 0.070 197.015 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.765 0.070 198.835 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.585 0.070 200.655 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.405 0.070 202.475 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.225 0.070 204.295 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.045 0.070 206.115 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.865 0.070 207.935 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.685 0.070 209.755 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.505 0.070 211.575 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.325 0.070 213.395 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.145 0.070 215.215 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.965 0.070 217.035 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.785 0.070 218.855 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.605 0.070 220.675 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.425 0.070 222.495 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.245 0.070 224.315 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.065 0.070 226.135 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.885 0.070 227.955 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.705 0.070 229.775 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.525 0.070 231.595 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.345 0.070 233.415 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.165 0.070 235.235 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.985 0.070 237.055 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.805 0.070 238.875 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.625 0.070 240.695 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.445 0.070 242.515 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.265 0.070 244.335 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.085 0.070 246.155 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.905 0.070 247.975 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.725 0.070 249.795 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.545 0.070 251.615 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.365 0.070 253.435 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.185 0.070 255.255 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.005 0.070 257.075 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.825 0.070 258.895 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.645 0.070 260.715 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.465 0.070 262.535 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.285 0.070 264.355 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.105 0.070 266.175 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.925 0.070 267.995 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.745 0.070 269.815 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.565 0.070 271.635 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.385 0.070 273.455 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.205 0.070 275.275 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.025 0.070 277.095 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.845 0.070 278.915 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.665 0.070 280.735 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.485 0.070 282.555 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.305 0.070 284.375 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.125 0.070 286.195 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.945 0.070 288.015 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.765 0.070 289.835 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.585 0.070 291.655 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.405 0.070 293.475 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.225 0.070 295.295 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.045 0.070 297.115 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.865 0.070 298.935 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.685 0.070 300.755 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.505 0.070 302.575 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.325 0.070 304.395 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.145 0.070 306.215 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.965 0.070 308.035 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.785 0.070 309.855 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.605 0.070 311.675 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.425 0.070 313.495 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.245 0.070 315.315 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.065 0.070 317.135 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.885 0.070 318.955 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.705 0.070 320.775 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.525 0.070 322.595 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.345 0.070 324.415 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.165 0.070 326.235 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.985 0.070 328.055 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.805 0.070 329.875 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.625 0.070 331.695 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.445 0.070 333.515 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.265 0.070 335.335 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.085 0.070 337.155 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.905 0.070 338.975 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.725 0.070 340.795 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.545 0.070 342.615 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.365 0.070 344.435 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.185 0.070 346.255 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.005 0.070 348.075 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.825 0.070 349.895 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.645 0.070 351.715 ;
    END
  END rd_out[95]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.125 0.070 356.195 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.945 0.070 358.015 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.765 0.070 359.835 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.585 0.070 361.655 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.405 0.070 363.475 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.225 0.070 365.295 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.045 0.070 367.115 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.865 0.070 368.935 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.685 0.070 370.755 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.505 0.070 372.575 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.325 0.070 374.395 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.145 0.070 376.215 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.965 0.070 378.035 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.785 0.070 379.855 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.605 0.070 381.675 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.425 0.070 383.495 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.245 0.070 385.315 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.065 0.070 387.135 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.885 0.070 388.955 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.705 0.070 390.775 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.525 0.070 392.595 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.345 0.070 394.415 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.165 0.070 396.235 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.985 0.070 398.055 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.805 0.070 399.875 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 401.625 0.070 401.695 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 403.445 0.070 403.515 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 405.265 0.070 405.335 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.085 0.070 407.155 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 408.905 0.070 408.975 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.725 0.070 410.795 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 412.545 0.070 412.615 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.365 0.070 414.435 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.185 0.070 416.255 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.005 0.070 418.075 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.825 0.070 419.895 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.645 0.070 421.715 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.465 0.070 423.535 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.285 0.070 425.355 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.105 0.070 427.175 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.925 0.070 428.995 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.745 0.070 430.815 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.565 0.070 432.635 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 434.385 0.070 434.455 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.205 0.070 436.275 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.025 0.070 438.095 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.845 0.070 439.915 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 441.665 0.070 441.735 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.485 0.070 443.555 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 445.305 0.070 445.375 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 447.125 0.070 447.195 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.945 0.070 449.015 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 450.765 0.070 450.835 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 452.585 0.070 452.655 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.405 0.070 454.475 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 456.225 0.070 456.295 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 458.045 0.070 458.115 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 459.865 0.070 459.935 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 461.685 0.070 461.755 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 463.505 0.070 463.575 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.325 0.070 465.395 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 467.145 0.070 467.215 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.965 0.070 469.035 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.785 0.070 470.855 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.605 0.070 472.675 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.425 0.070 474.495 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.245 0.070 476.315 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 478.065 0.070 478.135 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.885 0.070 479.955 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.705 0.070 481.775 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 483.525 0.070 483.595 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 485.345 0.070 485.415 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 487.165 0.070 487.235 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 488.985 0.070 489.055 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 490.805 0.070 490.875 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 492.625 0.070 492.695 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 494.445 0.070 494.515 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 496.265 0.070 496.335 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 498.085 0.070 498.155 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 499.905 0.070 499.975 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 501.725 0.070 501.795 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 503.545 0.070 503.615 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.365 0.070 505.435 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.185 0.070 507.255 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.005 0.070 509.075 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.825 0.070 510.895 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.645 0.070 512.715 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.465 0.070 514.535 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.285 0.070 516.355 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.105 0.070 518.175 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.925 0.070 519.995 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.745 0.070 521.815 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.565 0.070 523.635 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.385 0.070 525.455 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.205 0.070 527.275 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.025 0.070 529.095 ;
    END
  END wd_in[95]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.505 0.070 533.575 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.325 0.070 535.395 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.145 0.070 537.215 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.965 0.070 539.035 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.785 0.070 540.855 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.605 0.070 542.675 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.425 0.070 544.495 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.245 0.070 546.315 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.065 0.070 548.135 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.885 0.070 549.955 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.705 0.070 551.775 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.525 0.070 553.595 ;
    END
  END addr_in[11]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.005 0.070 558.075 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.825 0.070 559.895 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.645 0.070 561.715 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 571.200 ;
      RECT 3.500 1.400 3.780 571.200 ;
      RECT 5.740 1.400 6.020 571.200 ;
      RECT 7.980 1.400 8.260 571.200 ;
      RECT 10.220 1.400 10.500 571.200 ;
      RECT 12.460 1.400 12.740 571.200 ;
      RECT 14.700 1.400 14.980 571.200 ;
      RECT 16.940 1.400 17.220 571.200 ;
      RECT 19.180 1.400 19.460 571.200 ;
      RECT 21.420 1.400 21.700 571.200 ;
      RECT 23.660 1.400 23.940 571.200 ;
      RECT 25.900 1.400 26.180 571.200 ;
      RECT 28.140 1.400 28.420 571.200 ;
      RECT 30.380 1.400 30.660 571.200 ;
      RECT 32.620 1.400 32.900 571.200 ;
      RECT 34.860 1.400 35.140 571.200 ;
      RECT 37.100 1.400 37.380 571.200 ;
      RECT 39.340 1.400 39.620 571.200 ;
      RECT 41.580 1.400 41.860 571.200 ;
      RECT 43.820 1.400 44.100 571.200 ;
      RECT 46.060 1.400 46.340 571.200 ;
      RECT 48.300 1.400 48.580 571.200 ;
      RECT 50.540 1.400 50.820 571.200 ;
      RECT 52.780 1.400 53.060 571.200 ;
      RECT 55.020 1.400 55.300 571.200 ;
      RECT 57.260 1.400 57.540 571.200 ;
      RECT 59.500 1.400 59.780 571.200 ;
      RECT 61.740 1.400 62.020 571.200 ;
      RECT 63.980 1.400 64.260 571.200 ;
      RECT 66.220 1.400 66.500 571.200 ;
      RECT 68.460 1.400 68.740 571.200 ;
      RECT 70.700 1.400 70.980 571.200 ;
      RECT 72.940 1.400 73.220 571.200 ;
      RECT 75.180 1.400 75.460 571.200 ;
      RECT 77.420 1.400 77.700 571.200 ;
      RECT 79.660 1.400 79.940 571.200 ;
      RECT 81.900 1.400 82.180 571.200 ;
      RECT 84.140 1.400 84.420 571.200 ;
      RECT 86.380 1.400 86.660 571.200 ;
      RECT 88.620 1.400 88.900 571.200 ;
      RECT 90.860 1.400 91.140 571.200 ;
      RECT 93.100 1.400 93.380 571.200 ;
      RECT 95.340 1.400 95.620 571.200 ;
      RECT 97.580 1.400 97.860 571.200 ;
      RECT 99.820 1.400 100.100 571.200 ;
      RECT 102.060 1.400 102.340 571.200 ;
      RECT 104.300 1.400 104.580 571.200 ;
      RECT 106.540 1.400 106.820 571.200 ;
      RECT 108.780 1.400 109.060 571.200 ;
      RECT 111.020 1.400 111.300 571.200 ;
      RECT 113.260 1.400 113.540 571.200 ;
      RECT 115.500 1.400 115.780 571.200 ;
      RECT 117.740 1.400 118.020 571.200 ;
      RECT 119.980 1.400 120.260 571.200 ;
      RECT 122.220 1.400 122.500 571.200 ;
      RECT 124.460 1.400 124.740 571.200 ;
      RECT 126.700 1.400 126.980 571.200 ;
      RECT 128.940 1.400 129.220 571.200 ;
      RECT 131.180 1.400 131.460 571.200 ;
      RECT 133.420 1.400 133.700 571.200 ;
      RECT 135.660 1.400 135.940 571.200 ;
      RECT 137.900 1.400 138.180 571.200 ;
      RECT 140.140 1.400 140.420 571.200 ;
      RECT 142.380 1.400 142.660 571.200 ;
      RECT 144.620 1.400 144.900 571.200 ;
      RECT 146.860 1.400 147.140 571.200 ;
      RECT 149.100 1.400 149.380 571.200 ;
      RECT 151.340 1.400 151.620 571.200 ;
      RECT 153.580 1.400 153.860 571.200 ;
      RECT 155.820 1.400 156.100 571.200 ;
      RECT 158.060 1.400 158.340 571.200 ;
      RECT 160.300 1.400 160.580 571.200 ;
      RECT 162.540 1.400 162.820 571.200 ;
      RECT 164.780 1.400 165.060 571.200 ;
      RECT 167.020 1.400 167.300 571.200 ;
      RECT 169.260 1.400 169.540 571.200 ;
      RECT 171.500 1.400 171.780 571.200 ;
      RECT 173.740 1.400 174.020 571.200 ;
      RECT 175.980 1.400 176.260 571.200 ;
      RECT 178.220 1.400 178.500 571.200 ;
      RECT 180.460 1.400 180.740 571.200 ;
      RECT 182.700 1.400 182.980 571.200 ;
      RECT 184.940 1.400 185.220 571.200 ;
      RECT 187.180 1.400 187.460 571.200 ;
      RECT 189.420 1.400 189.700 571.200 ;
      RECT 191.660 1.400 191.940 571.200 ;
      RECT 193.900 1.400 194.180 571.200 ;
      RECT 196.140 1.400 196.420 571.200 ;
      RECT 198.380 1.400 198.660 571.200 ;
      RECT 200.620 1.400 200.900 571.200 ;
      RECT 202.860 1.400 203.140 571.200 ;
      RECT 205.100 1.400 205.380 571.200 ;
      RECT 207.340 1.400 207.620 571.200 ;
      RECT 209.580 1.400 209.860 571.200 ;
      RECT 211.820 1.400 212.100 571.200 ;
      RECT 214.060 1.400 214.340 571.200 ;
      RECT 216.300 1.400 216.580 571.200 ;
      RECT 218.540 1.400 218.820 571.200 ;
      RECT 220.780 1.400 221.060 571.200 ;
      RECT 223.020 1.400 223.300 571.200 ;
      RECT 225.260 1.400 225.540 571.200 ;
      RECT 227.500 1.400 227.780 571.200 ;
      RECT 229.740 1.400 230.020 571.200 ;
      RECT 231.980 1.400 232.260 571.200 ;
      RECT 234.220 1.400 234.500 571.200 ;
      RECT 236.460 1.400 236.740 571.200 ;
      RECT 238.700 1.400 238.980 571.200 ;
      RECT 240.940 1.400 241.220 571.200 ;
      RECT 243.180 1.400 243.460 571.200 ;
      RECT 245.420 1.400 245.700 571.200 ;
      RECT 247.660 1.400 247.940 571.200 ;
      RECT 249.900 1.400 250.180 571.200 ;
      RECT 252.140 1.400 252.420 571.200 ;
      RECT 254.380 1.400 254.660 571.200 ;
      RECT 256.620 1.400 256.900 571.200 ;
      RECT 258.860 1.400 259.140 571.200 ;
      RECT 261.100 1.400 261.380 571.200 ;
      RECT 263.340 1.400 263.620 571.200 ;
      RECT 265.580 1.400 265.860 571.200 ;
      RECT 267.820 1.400 268.100 571.200 ;
      RECT 270.060 1.400 270.340 571.200 ;
      RECT 272.300 1.400 272.580 571.200 ;
      RECT 274.540 1.400 274.820 571.200 ;
      RECT 276.780 1.400 277.060 571.200 ;
      RECT 279.020 1.400 279.300 571.200 ;
      RECT 281.260 1.400 281.540 571.200 ;
      RECT 283.500 1.400 283.780 571.200 ;
      RECT 285.740 1.400 286.020 571.200 ;
      RECT 287.980 1.400 288.260 571.200 ;
      RECT 290.220 1.400 290.500 571.200 ;
      RECT 292.460 1.400 292.740 571.200 ;
      RECT 294.700 1.400 294.980 571.200 ;
      RECT 296.940 1.400 297.220 571.200 ;
      RECT 299.180 1.400 299.460 571.200 ;
      RECT 301.420 1.400 301.700 571.200 ;
      RECT 303.660 1.400 303.940 571.200 ;
      RECT 305.900 1.400 306.180 571.200 ;
      RECT 308.140 1.400 308.420 571.200 ;
      RECT 310.380 1.400 310.660 571.200 ;
      RECT 312.620 1.400 312.900 571.200 ;
      RECT 314.860 1.400 315.140 571.200 ;
      RECT 317.100 1.400 317.380 571.200 ;
      RECT 319.340 1.400 319.620 571.200 ;
      RECT 321.580 1.400 321.860 571.200 ;
      RECT 323.820 1.400 324.100 571.200 ;
      RECT 326.060 1.400 326.340 571.200 ;
      RECT 328.300 1.400 328.580 571.200 ;
      RECT 330.540 1.400 330.820 571.200 ;
      RECT 332.780 1.400 333.060 571.200 ;
      RECT 335.020 1.400 335.300 571.200 ;
      RECT 337.260 1.400 337.540 571.200 ;
      RECT 339.500 1.400 339.780 571.200 ;
      RECT 341.740 1.400 342.020 571.200 ;
      RECT 343.980 1.400 344.260 571.200 ;
      RECT 346.220 1.400 346.500 571.200 ;
      RECT 348.460 1.400 348.740 571.200 ;
      RECT 350.700 1.400 350.980 571.200 ;
      RECT 352.940 1.400 353.220 571.200 ;
      RECT 355.180 1.400 355.460 571.200 ;
      RECT 357.420 1.400 357.700 571.200 ;
      RECT 359.660 1.400 359.940 571.200 ;
      RECT 361.900 1.400 362.180 571.200 ;
      RECT 364.140 1.400 364.420 571.200 ;
      RECT 366.380 1.400 366.660 571.200 ;
      RECT 368.620 1.400 368.900 571.200 ;
      RECT 370.860 1.400 371.140 571.200 ;
      RECT 373.100 1.400 373.380 571.200 ;
      RECT 375.340 1.400 375.620 571.200 ;
      RECT 377.580 1.400 377.860 571.200 ;
      RECT 379.820 1.400 380.100 571.200 ;
      RECT 382.060 1.400 382.340 571.200 ;
      RECT 384.300 1.400 384.580 571.200 ;
      RECT 386.540 1.400 386.820 571.200 ;
      RECT 388.780 1.400 389.060 571.200 ;
      RECT 391.020 1.400 391.300 571.200 ;
      RECT 393.260 1.400 393.540 571.200 ;
      RECT 395.500 1.400 395.780 571.200 ;
      RECT 397.740 1.400 398.020 571.200 ;
      RECT 399.980 1.400 400.260 571.200 ;
      RECT 402.220 1.400 402.500 571.200 ;
      RECT 404.460 1.400 404.740 571.200 ;
      RECT 406.700 1.400 406.980 571.200 ;
      RECT 408.940 1.400 409.220 571.200 ;
      RECT 411.180 1.400 411.460 571.200 ;
      RECT 413.420 1.400 413.700 571.200 ;
      RECT 415.660 1.400 415.940 571.200 ;
      RECT 417.900 1.400 418.180 571.200 ;
      RECT 420.140 1.400 420.420 571.200 ;
      RECT 422.380 1.400 422.660 571.200 ;
      RECT 424.620 1.400 424.900 571.200 ;
      RECT 426.860 1.400 427.140 571.200 ;
      RECT 429.100 1.400 429.380 571.200 ;
      RECT 431.340 1.400 431.620 571.200 ;
      RECT 433.580 1.400 433.860 571.200 ;
      RECT 435.820 1.400 436.100 571.200 ;
      RECT 438.060 1.400 438.340 571.200 ;
      RECT 440.300 1.400 440.580 571.200 ;
      RECT 442.540 1.400 442.820 571.200 ;
      RECT 444.780 1.400 445.060 571.200 ;
      RECT 447.020 1.400 447.300 571.200 ;
      RECT 449.260 1.400 449.540 571.200 ;
      RECT 451.500 1.400 451.780 571.200 ;
      RECT 453.740 1.400 454.020 571.200 ;
      RECT 455.980 1.400 456.260 571.200 ;
      RECT 458.220 1.400 458.500 571.200 ;
      RECT 460.460 1.400 460.740 571.200 ;
      RECT 462.700 1.400 462.980 571.200 ;
      RECT 464.940 1.400 465.220 571.200 ;
      RECT 467.180 1.400 467.460 571.200 ;
      RECT 469.420 1.400 469.700 571.200 ;
      RECT 471.660 1.400 471.940 571.200 ;
      RECT 473.900 1.400 474.180 571.200 ;
      RECT 476.140 1.400 476.420 571.200 ;
      RECT 478.380 1.400 478.660 571.200 ;
      RECT 480.620 1.400 480.900 571.200 ;
      RECT 482.860 1.400 483.140 571.200 ;
      RECT 485.100 1.400 485.380 571.200 ;
      RECT 487.340 1.400 487.620 571.200 ;
      RECT 489.580 1.400 489.860 571.200 ;
      RECT 491.820 1.400 492.100 571.200 ;
      RECT 494.060 1.400 494.340 571.200 ;
      RECT 496.300 1.400 496.580 571.200 ;
      RECT 498.540 1.400 498.820 571.200 ;
      RECT 500.780 1.400 501.060 571.200 ;
      RECT 503.020 1.400 503.300 571.200 ;
      RECT 505.260 1.400 505.540 571.200 ;
      RECT 507.500 1.400 507.780 571.200 ;
      RECT 509.740 1.400 510.020 571.200 ;
      RECT 511.980 1.400 512.260 571.200 ;
      RECT 514.220 1.400 514.500 571.200 ;
      RECT 516.460 1.400 516.740 571.200 ;
      RECT 518.700 1.400 518.980 571.200 ;
      RECT 520.940 1.400 521.220 571.200 ;
      RECT 523.180 1.400 523.460 571.200 ;
      RECT 525.420 1.400 525.700 571.200 ;
      RECT 527.660 1.400 527.940 571.200 ;
      RECT 529.900 1.400 530.180 571.200 ;
      RECT 532.140 1.400 532.420 571.200 ;
      RECT 534.380 1.400 534.660 571.200 ;
      RECT 536.620 1.400 536.900 571.200 ;
      RECT 538.860 1.400 539.140 571.200 ;
      RECT 541.100 1.400 541.380 571.200 ;
      RECT 543.340 1.400 543.620 571.200 ;
      RECT 545.580 1.400 545.860 571.200 ;
      RECT 547.820 1.400 548.100 571.200 ;
      RECT 550.060 1.400 550.340 571.200 ;
      RECT 552.300 1.400 552.580 571.200 ;
      RECT 554.540 1.400 554.820 571.200 ;
      RECT 556.780 1.400 557.060 571.200 ;
      RECT 559.020 1.400 559.300 571.200 ;
      RECT 561.260 1.400 561.540 571.200 ;
      RECT 563.500 1.400 563.780 571.200 ;
      RECT 565.740 1.400 566.020 571.200 ;
      RECT 567.980 1.400 568.260 571.200 ;
      RECT 570.220 1.400 570.500 571.200 ;
      RECT 572.460 1.400 572.740 571.200 ;
      RECT 574.700 1.400 574.980 571.200 ;
      RECT 576.940 1.400 577.220 571.200 ;
      RECT 579.180 1.400 579.460 571.200 ;
      RECT 581.420 1.400 581.700 571.200 ;
      RECT 583.660 1.400 583.940 571.200 ;
      RECT 585.900 1.400 586.180 571.200 ;
      RECT 588.140 1.400 588.420 571.200 ;
      RECT 590.380 1.400 590.660 571.200 ;
      RECT 592.620 1.400 592.900 571.200 ;
      RECT 594.860 1.400 595.140 571.200 ;
      RECT 597.100 1.400 597.380 571.200 ;
      RECT 599.340 1.400 599.620 571.200 ;
      RECT 601.580 1.400 601.860 571.200 ;
      RECT 603.820 1.400 604.100 571.200 ;
      RECT 606.060 1.400 606.340 571.200 ;
      RECT 608.300 1.400 608.580 571.200 ;
      RECT 610.540 1.400 610.820 571.200 ;
      RECT 612.780 1.400 613.060 571.200 ;
      RECT 615.020 1.400 615.300 571.200 ;
      RECT 617.260 1.400 617.540 571.200 ;
      RECT 619.500 1.400 619.780 571.200 ;
      RECT 621.740 1.400 622.020 571.200 ;
      RECT 623.980 1.400 624.260 571.200 ;
      RECT 626.220 1.400 626.500 571.200 ;
      RECT 628.460 1.400 628.740 571.200 ;
      RECT 630.700 1.400 630.980 571.200 ;
      RECT 632.940 1.400 633.220 571.200 ;
      RECT 635.180 1.400 635.460 571.200 ;
      RECT 637.420 1.400 637.700 571.200 ;
      RECT 639.660 1.400 639.940 571.200 ;
      RECT 641.900 1.400 642.180 571.200 ;
      RECT 644.140 1.400 644.420 571.200 ;
      RECT 646.380 1.400 646.660 571.200 ;
      RECT 648.620 1.400 648.900 571.200 ;
      RECT 650.860 1.400 651.140 571.200 ;
      RECT 653.100 1.400 653.380 571.200 ;
      RECT 655.340 1.400 655.620 571.200 ;
      RECT 657.580 1.400 657.860 571.200 ;
      RECT 659.820 1.400 660.100 571.200 ;
      RECT 662.060 1.400 662.340 571.200 ;
      RECT 664.300 1.400 664.580 571.200 ;
      RECT 666.540 1.400 666.820 571.200 ;
      RECT 668.780 1.400 669.060 571.200 ;
      RECT 671.020 1.400 671.300 571.200 ;
      RECT 673.260 1.400 673.540 571.200 ;
      RECT 675.500 1.400 675.780 571.200 ;
      RECT 677.740 1.400 678.020 571.200 ;
      RECT 679.980 1.400 680.260 571.200 ;
      RECT 682.220 1.400 682.500 571.200 ;
      RECT 684.460 1.400 684.740 571.200 ;
      RECT 686.700 1.400 686.980 571.200 ;
      RECT 688.940 1.400 689.220 571.200 ;
      RECT 691.180 1.400 691.460 571.200 ;
      RECT 693.420 1.400 693.700 571.200 ;
      RECT 695.660 1.400 695.940 571.200 ;
      RECT 697.900 1.400 698.180 571.200 ;
      RECT 700.140 1.400 700.420 571.200 ;
      RECT 702.380 1.400 702.660 571.200 ;
      RECT 704.620 1.400 704.900 571.200 ;
      RECT 706.860 1.400 707.140 571.200 ;
      RECT 709.100 1.400 709.380 571.200 ;
      RECT 711.340 1.400 711.620 571.200 ;
      RECT 713.580 1.400 713.860 571.200 ;
      RECT 715.820 1.400 716.100 571.200 ;
      RECT 718.060 1.400 718.340 571.200 ;
      RECT 720.300 1.400 720.580 571.200 ;
      RECT 722.540 1.400 722.820 571.200 ;
      RECT 724.780 1.400 725.060 571.200 ;
      RECT 727.020 1.400 727.300 571.200 ;
      RECT 729.260 1.400 729.540 571.200 ;
      RECT 731.500 1.400 731.780 571.200 ;
      RECT 733.740 1.400 734.020 571.200 ;
      RECT 735.980 1.400 736.260 571.200 ;
      RECT 738.220 1.400 738.500 571.200 ;
      RECT 740.460 1.400 740.740 571.200 ;
      RECT 742.700 1.400 742.980 571.200 ;
      RECT 744.940 1.400 745.220 571.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 571.200 ;
      RECT 4.620 1.400 4.900 571.200 ;
      RECT 6.860 1.400 7.140 571.200 ;
      RECT 9.100 1.400 9.380 571.200 ;
      RECT 11.340 1.400 11.620 571.200 ;
      RECT 13.580 1.400 13.860 571.200 ;
      RECT 15.820 1.400 16.100 571.200 ;
      RECT 18.060 1.400 18.340 571.200 ;
      RECT 20.300 1.400 20.580 571.200 ;
      RECT 22.540 1.400 22.820 571.200 ;
      RECT 24.780 1.400 25.060 571.200 ;
      RECT 27.020 1.400 27.300 571.200 ;
      RECT 29.260 1.400 29.540 571.200 ;
      RECT 31.500 1.400 31.780 571.200 ;
      RECT 33.740 1.400 34.020 571.200 ;
      RECT 35.980 1.400 36.260 571.200 ;
      RECT 38.220 1.400 38.500 571.200 ;
      RECT 40.460 1.400 40.740 571.200 ;
      RECT 42.700 1.400 42.980 571.200 ;
      RECT 44.940 1.400 45.220 571.200 ;
      RECT 47.180 1.400 47.460 571.200 ;
      RECT 49.420 1.400 49.700 571.200 ;
      RECT 51.660 1.400 51.940 571.200 ;
      RECT 53.900 1.400 54.180 571.200 ;
      RECT 56.140 1.400 56.420 571.200 ;
      RECT 58.380 1.400 58.660 571.200 ;
      RECT 60.620 1.400 60.900 571.200 ;
      RECT 62.860 1.400 63.140 571.200 ;
      RECT 65.100 1.400 65.380 571.200 ;
      RECT 67.340 1.400 67.620 571.200 ;
      RECT 69.580 1.400 69.860 571.200 ;
      RECT 71.820 1.400 72.100 571.200 ;
      RECT 74.060 1.400 74.340 571.200 ;
      RECT 76.300 1.400 76.580 571.200 ;
      RECT 78.540 1.400 78.820 571.200 ;
      RECT 80.780 1.400 81.060 571.200 ;
      RECT 83.020 1.400 83.300 571.200 ;
      RECT 85.260 1.400 85.540 571.200 ;
      RECT 87.500 1.400 87.780 571.200 ;
      RECT 89.740 1.400 90.020 571.200 ;
      RECT 91.980 1.400 92.260 571.200 ;
      RECT 94.220 1.400 94.500 571.200 ;
      RECT 96.460 1.400 96.740 571.200 ;
      RECT 98.700 1.400 98.980 571.200 ;
      RECT 100.940 1.400 101.220 571.200 ;
      RECT 103.180 1.400 103.460 571.200 ;
      RECT 105.420 1.400 105.700 571.200 ;
      RECT 107.660 1.400 107.940 571.200 ;
      RECT 109.900 1.400 110.180 571.200 ;
      RECT 112.140 1.400 112.420 571.200 ;
      RECT 114.380 1.400 114.660 571.200 ;
      RECT 116.620 1.400 116.900 571.200 ;
      RECT 118.860 1.400 119.140 571.200 ;
      RECT 121.100 1.400 121.380 571.200 ;
      RECT 123.340 1.400 123.620 571.200 ;
      RECT 125.580 1.400 125.860 571.200 ;
      RECT 127.820 1.400 128.100 571.200 ;
      RECT 130.060 1.400 130.340 571.200 ;
      RECT 132.300 1.400 132.580 571.200 ;
      RECT 134.540 1.400 134.820 571.200 ;
      RECT 136.780 1.400 137.060 571.200 ;
      RECT 139.020 1.400 139.300 571.200 ;
      RECT 141.260 1.400 141.540 571.200 ;
      RECT 143.500 1.400 143.780 571.200 ;
      RECT 145.740 1.400 146.020 571.200 ;
      RECT 147.980 1.400 148.260 571.200 ;
      RECT 150.220 1.400 150.500 571.200 ;
      RECT 152.460 1.400 152.740 571.200 ;
      RECT 154.700 1.400 154.980 571.200 ;
      RECT 156.940 1.400 157.220 571.200 ;
      RECT 159.180 1.400 159.460 571.200 ;
      RECT 161.420 1.400 161.700 571.200 ;
      RECT 163.660 1.400 163.940 571.200 ;
      RECT 165.900 1.400 166.180 571.200 ;
      RECT 168.140 1.400 168.420 571.200 ;
      RECT 170.380 1.400 170.660 571.200 ;
      RECT 172.620 1.400 172.900 571.200 ;
      RECT 174.860 1.400 175.140 571.200 ;
      RECT 177.100 1.400 177.380 571.200 ;
      RECT 179.340 1.400 179.620 571.200 ;
      RECT 181.580 1.400 181.860 571.200 ;
      RECT 183.820 1.400 184.100 571.200 ;
      RECT 186.060 1.400 186.340 571.200 ;
      RECT 188.300 1.400 188.580 571.200 ;
      RECT 190.540 1.400 190.820 571.200 ;
      RECT 192.780 1.400 193.060 571.200 ;
      RECT 195.020 1.400 195.300 571.200 ;
      RECT 197.260 1.400 197.540 571.200 ;
      RECT 199.500 1.400 199.780 571.200 ;
      RECT 201.740 1.400 202.020 571.200 ;
      RECT 203.980 1.400 204.260 571.200 ;
      RECT 206.220 1.400 206.500 571.200 ;
      RECT 208.460 1.400 208.740 571.200 ;
      RECT 210.700 1.400 210.980 571.200 ;
      RECT 212.940 1.400 213.220 571.200 ;
      RECT 215.180 1.400 215.460 571.200 ;
      RECT 217.420 1.400 217.700 571.200 ;
      RECT 219.660 1.400 219.940 571.200 ;
      RECT 221.900 1.400 222.180 571.200 ;
      RECT 224.140 1.400 224.420 571.200 ;
      RECT 226.380 1.400 226.660 571.200 ;
      RECT 228.620 1.400 228.900 571.200 ;
      RECT 230.860 1.400 231.140 571.200 ;
      RECT 233.100 1.400 233.380 571.200 ;
      RECT 235.340 1.400 235.620 571.200 ;
      RECT 237.580 1.400 237.860 571.200 ;
      RECT 239.820 1.400 240.100 571.200 ;
      RECT 242.060 1.400 242.340 571.200 ;
      RECT 244.300 1.400 244.580 571.200 ;
      RECT 246.540 1.400 246.820 571.200 ;
      RECT 248.780 1.400 249.060 571.200 ;
      RECT 251.020 1.400 251.300 571.200 ;
      RECT 253.260 1.400 253.540 571.200 ;
      RECT 255.500 1.400 255.780 571.200 ;
      RECT 257.740 1.400 258.020 571.200 ;
      RECT 259.980 1.400 260.260 571.200 ;
      RECT 262.220 1.400 262.500 571.200 ;
      RECT 264.460 1.400 264.740 571.200 ;
      RECT 266.700 1.400 266.980 571.200 ;
      RECT 268.940 1.400 269.220 571.200 ;
      RECT 271.180 1.400 271.460 571.200 ;
      RECT 273.420 1.400 273.700 571.200 ;
      RECT 275.660 1.400 275.940 571.200 ;
      RECT 277.900 1.400 278.180 571.200 ;
      RECT 280.140 1.400 280.420 571.200 ;
      RECT 282.380 1.400 282.660 571.200 ;
      RECT 284.620 1.400 284.900 571.200 ;
      RECT 286.860 1.400 287.140 571.200 ;
      RECT 289.100 1.400 289.380 571.200 ;
      RECT 291.340 1.400 291.620 571.200 ;
      RECT 293.580 1.400 293.860 571.200 ;
      RECT 295.820 1.400 296.100 571.200 ;
      RECT 298.060 1.400 298.340 571.200 ;
      RECT 300.300 1.400 300.580 571.200 ;
      RECT 302.540 1.400 302.820 571.200 ;
      RECT 304.780 1.400 305.060 571.200 ;
      RECT 307.020 1.400 307.300 571.200 ;
      RECT 309.260 1.400 309.540 571.200 ;
      RECT 311.500 1.400 311.780 571.200 ;
      RECT 313.740 1.400 314.020 571.200 ;
      RECT 315.980 1.400 316.260 571.200 ;
      RECT 318.220 1.400 318.500 571.200 ;
      RECT 320.460 1.400 320.740 571.200 ;
      RECT 322.700 1.400 322.980 571.200 ;
      RECT 324.940 1.400 325.220 571.200 ;
      RECT 327.180 1.400 327.460 571.200 ;
      RECT 329.420 1.400 329.700 571.200 ;
      RECT 331.660 1.400 331.940 571.200 ;
      RECT 333.900 1.400 334.180 571.200 ;
      RECT 336.140 1.400 336.420 571.200 ;
      RECT 338.380 1.400 338.660 571.200 ;
      RECT 340.620 1.400 340.900 571.200 ;
      RECT 342.860 1.400 343.140 571.200 ;
      RECT 345.100 1.400 345.380 571.200 ;
      RECT 347.340 1.400 347.620 571.200 ;
      RECT 349.580 1.400 349.860 571.200 ;
      RECT 351.820 1.400 352.100 571.200 ;
      RECT 354.060 1.400 354.340 571.200 ;
      RECT 356.300 1.400 356.580 571.200 ;
      RECT 358.540 1.400 358.820 571.200 ;
      RECT 360.780 1.400 361.060 571.200 ;
      RECT 363.020 1.400 363.300 571.200 ;
      RECT 365.260 1.400 365.540 571.200 ;
      RECT 367.500 1.400 367.780 571.200 ;
      RECT 369.740 1.400 370.020 571.200 ;
      RECT 371.980 1.400 372.260 571.200 ;
      RECT 374.220 1.400 374.500 571.200 ;
      RECT 376.460 1.400 376.740 571.200 ;
      RECT 378.700 1.400 378.980 571.200 ;
      RECT 380.940 1.400 381.220 571.200 ;
      RECT 383.180 1.400 383.460 571.200 ;
      RECT 385.420 1.400 385.700 571.200 ;
      RECT 387.660 1.400 387.940 571.200 ;
      RECT 389.900 1.400 390.180 571.200 ;
      RECT 392.140 1.400 392.420 571.200 ;
      RECT 394.380 1.400 394.660 571.200 ;
      RECT 396.620 1.400 396.900 571.200 ;
      RECT 398.860 1.400 399.140 571.200 ;
      RECT 401.100 1.400 401.380 571.200 ;
      RECT 403.340 1.400 403.620 571.200 ;
      RECT 405.580 1.400 405.860 571.200 ;
      RECT 407.820 1.400 408.100 571.200 ;
      RECT 410.060 1.400 410.340 571.200 ;
      RECT 412.300 1.400 412.580 571.200 ;
      RECT 414.540 1.400 414.820 571.200 ;
      RECT 416.780 1.400 417.060 571.200 ;
      RECT 419.020 1.400 419.300 571.200 ;
      RECT 421.260 1.400 421.540 571.200 ;
      RECT 423.500 1.400 423.780 571.200 ;
      RECT 425.740 1.400 426.020 571.200 ;
      RECT 427.980 1.400 428.260 571.200 ;
      RECT 430.220 1.400 430.500 571.200 ;
      RECT 432.460 1.400 432.740 571.200 ;
      RECT 434.700 1.400 434.980 571.200 ;
      RECT 436.940 1.400 437.220 571.200 ;
      RECT 439.180 1.400 439.460 571.200 ;
      RECT 441.420 1.400 441.700 571.200 ;
      RECT 443.660 1.400 443.940 571.200 ;
      RECT 445.900 1.400 446.180 571.200 ;
      RECT 448.140 1.400 448.420 571.200 ;
      RECT 450.380 1.400 450.660 571.200 ;
      RECT 452.620 1.400 452.900 571.200 ;
      RECT 454.860 1.400 455.140 571.200 ;
      RECT 457.100 1.400 457.380 571.200 ;
      RECT 459.340 1.400 459.620 571.200 ;
      RECT 461.580 1.400 461.860 571.200 ;
      RECT 463.820 1.400 464.100 571.200 ;
      RECT 466.060 1.400 466.340 571.200 ;
      RECT 468.300 1.400 468.580 571.200 ;
      RECT 470.540 1.400 470.820 571.200 ;
      RECT 472.780 1.400 473.060 571.200 ;
      RECT 475.020 1.400 475.300 571.200 ;
      RECT 477.260 1.400 477.540 571.200 ;
      RECT 479.500 1.400 479.780 571.200 ;
      RECT 481.740 1.400 482.020 571.200 ;
      RECT 483.980 1.400 484.260 571.200 ;
      RECT 486.220 1.400 486.500 571.200 ;
      RECT 488.460 1.400 488.740 571.200 ;
      RECT 490.700 1.400 490.980 571.200 ;
      RECT 492.940 1.400 493.220 571.200 ;
      RECT 495.180 1.400 495.460 571.200 ;
      RECT 497.420 1.400 497.700 571.200 ;
      RECT 499.660 1.400 499.940 571.200 ;
      RECT 501.900 1.400 502.180 571.200 ;
      RECT 504.140 1.400 504.420 571.200 ;
      RECT 506.380 1.400 506.660 571.200 ;
      RECT 508.620 1.400 508.900 571.200 ;
      RECT 510.860 1.400 511.140 571.200 ;
      RECT 513.100 1.400 513.380 571.200 ;
      RECT 515.340 1.400 515.620 571.200 ;
      RECT 517.580 1.400 517.860 571.200 ;
      RECT 519.820 1.400 520.100 571.200 ;
      RECT 522.060 1.400 522.340 571.200 ;
      RECT 524.300 1.400 524.580 571.200 ;
      RECT 526.540 1.400 526.820 571.200 ;
      RECT 528.780 1.400 529.060 571.200 ;
      RECT 531.020 1.400 531.300 571.200 ;
      RECT 533.260 1.400 533.540 571.200 ;
      RECT 535.500 1.400 535.780 571.200 ;
      RECT 537.740 1.400 538.020 571.200 ;
      RECT 539.980 1.400 540.260 571.200 ;
      RECT 542.220 1.400 542.500 571.200 ;
      RECT 544.460 1.400 544.740 571.200 ;
      RECT 546.700 1.400 546.980 571.200 ;
      RECT 548.940 1.400 549.220 571.200 ;
      RECT 551.180 1.400 551.460 571.200 ;
      RECT 553.420 1.400 553.700 571.200 ;
      RECT 555.660 1.400 555.940 571.200 ;
      RECT 557.900 1.400 558.180 571.200 ;
      RECT 560.140 1.400 560.420 571.200 ;
      RECT 562.380 1.400 562.660 571.200 ;
      RECT 564.620 1.400 564.900 571.200 ;
      RECT 566.860 1.400 567.140 571.200 ;
      RECT 569.100 1.400 569.380 571.200 ;
      RECT 571.340 1.400 571.620 571.200 ;
      RECT 573.580 1.400 573.860 571.200 ;
      RECT 575.820 1.400 576.100 571.200 ;
      RECT 578.060 1.400 578.340 571.200 ;
      RECT 580.300 1.400 580.580 571.200 ;
      RECT 582.540 1.400 582.820 571.200 ;
      RECT 584.780 1.400 585.060 571.200 ;
      RECT 587.020 1.400 587.300 571.200 ;
      RECT 589.260 1.400 589.540 571.200 ;
      RECT 591.500 1.400 591.780 571.200 ;
      RECT 593.740 1.400 594.020 571.200 ;
      RECT 595.980 1.400 596.260 571.200 ;
      RECT 598.220 1.400 598.500 571.200 ;
      RECT 600.460 1.400 600.740 571.200 ;
      RECT 602.700 1.400 602.980 571.200 ;
      RECT 604.940 1.400 605.220 571.200 ;
      RECT 607.180 1.400 607.460 571.200 ;
      RECT 609.420 1.400 609.700 571.200 ;
      RECT 611.660 1.400 611.940 571.200 ;
      RECT 613.900 1.400 614.180 571.200 ;
      RECT 616.140 1.400 616.420 571.200 ;
      RECT 618.380 1.400 618.660 571.200 ;
      RECT 620.620 1.400 620.900 571.200 ;
      RECT 622.860 1.400 623.140 571.200 ;
      RECT 625.100 1.400 625.380 571.200 ;
      RECT 627.340 1.400 627.620 571.200 ;
      RECT 629.580 1.400 629.860 571.200 ;
      RECT 631.820 1.400 632.100 571.200 ;
      RECT 634.060 1.400 634.340 571.200 ;
      RECT 636.300 1.400 636.580 571.200 ;
      RECT 638.540 1.400 638.820 571.200 ;
      RECT 640.780 1.400 641.060 571.200 ;
      RECT 643.020 1.400 643.300 571.200 ;
      RECT 645.260 1.400 645.540 571.200 ;
      RECT 647.500 1.400 647.780 571.200 ;
      RECT 649.740 1.400 650.020 571.200 ;
      RECT 651.980 1.400 652.260 571.200 ;
      RECT 654.220 1.400 654.500 571.200 ;
      RECT 656.460 1.400 656.740 571.200 ;
      RECT 658.700 1.400 658.980 571.200 ;
      RECT 660.940 1.400 661.220 571.200 ;
      RECT 663.180 1.400 663.460 571.200 ;
      RECT 665.420 1.400 665.700 571.200 ;
      RECT 667.660 1.400 667.940 571.200 ;
      RECT 669.900 1.400 670.180 571.200 ;
      RECT 672.140 1.400 672.420 571.200 ;
      RECT 674.380 1.400 674.660 571.200 ;
      RECT 676.620 1.400 676.900 571.200 ;
      RECT 678.860 1.400 679.140 571.200 ;
      RECT 681.100 1.400 681.380 571.200 ;
      RECT 683.340 1.400 683.620 571.200 ;
      RECT 685.580 1.400 685.860 571.200 ;
      RECT 687.820 1.400 688.100 571.200 ;
      RECT 690.060 1.400 690.340 571.200 ;
      RECT 692.300 1.400 692.580 571.200 ;
      RECT 694.540 1.400 694.820 571.200 ;
      RECT 696.780 1.400 697.060 571.200 ;
      RECT 699.020 1.400 699.300 571.200 ;
      RECT 701.260 1.400 701.540 571.200 ;
      RECT 703.500 1.400 703.780 571.200 ;
      RECT 705.740 1.400 706.020 571.200 ;
      RECT 707.980 1.400 708.260 571.200 ;
      RECT 710.220 1.400 710.500 571.200 ;
      RECT 712.460 1.400 712.740 571.200 ;
      RECT 714.700 1.400 714.980 571.200 ;
      RECT 716.940 1.400 717.220 571.200 ;
      RECT 719.180 1.400 719.460 571.200 ;
      RECT 721.420 1.400 721.700 571.200 ;
      RECT 723.660 1.400 723.940 571.200 ;
      RECT 725.900 1.400 726.180 571.200 ;
      RECT 728.140 1.400 728.420 571.200 ;
      RECT 730.380 1.400 730.660 571.200 ;
      RECT 732.620 1.400 732.900 571.200 ;
      RECT 734.860 1.400 735.140 571.200 ;
      RECT 737.100 1.400 737.380 571.200 ;
      RECT 739.340 1.400 739.620 571.200 ;
      RECT 741.580 1.400 741.860 571.200 ;
      RECT 743.820 1.400 744.100 571.200 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 747.080 572.600 ;
    LAYER metal2 ;
    RECT 0 0 747.080 572.600 ;
    LAYER metal3 ;
    RECT 0.070 0 747.080 572.600 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 3.185 ;
    RECT 0 3.255 0.070 5.005 ;
    RECT 0 5.075 0.070 6.825 ;
    RECT 0 6.895 0.070 8.645 ;
    RECT 0 8.715 0.070 10.465 ;
    RECT 0 10.535 0.070 12.285 ;
    RECT 0 12.355 0.070 14.105 ;
    RECT 0 14.175 0.070 15.925 ;
    RECT 0 15.995 0.070 17.745 ;
    RECT 0 17.815 0.070 19.565 ;
    RECT 0 19.635 0.070 21.385 ;
    RECT 0 21.455 0.070 23.205 ;
    RECT 0 23.275 0.070 25.025 ;
    RECT 0 25.095 0.070 26.845 ;
    RECT 0 26.915 0.070 28.665 ;
    RECT 0 28.735 0.070 30.485 ;
    RECT 0 30.555 0.070 32.305 ;
    RECT 0 32.375 0.070 34.125 ;
    RECT 0 34.195 0.070 35.945 ;
    RECT 0 36.015 0.070 37.765 ;
    RECT 0 37.835 0.070 39.585 ;
    RECT 0 39.655 0.070 41.405 ;
    RECT 0 41.475 0.070 43.225 ;
    RECT 0 43.295 0.070 45.045 ;
    RECT 0 45.115 0.070 46.865 ;
    RECT 0 46.935 0.070 48.685 ;
    RECT 0 48.755 0.070 50.505 ;
    RECT 0 50.575 0.070 52.325 ;
    RECT 0 52.395 0.070 54.145 ;
    RECT 0 54.215 0.070 55.965 ;
    RECT 0 56.035 0.070 57.785 ;
    RECT 0 57.855 0.070 59.605 ;
    RECT 0 59.675 0.070 61.425 ;
    RECT 0 61.495 0.070 63.245 ;
    RECT 0 63.315 0.070 65.065 ;
    RECT 0 65.135 0.070 66.885 ;
    RECT 0 66.955 0.070 68.705 ;
    RECT 0 68.775 0.070 70.525 ;
    RECT 0 70.595 0.070 72.345 ;
    RECT 0 72.415 0.070 74.165 ;
    RECT 0 74.235 0.070 75.985 ;
    RECT 0 76.055 0.070 77.805 ;
    RECT 0 77.875 0.070 79.625 ;
    RECT 0 79.695 0.070 81.445 ;
    RECT 0 81.515 0.070 83.265 ;
    RECT 0 83.335 0.070 85.085 ;
    RECT 0 85.155 0.070 86.905 ;
    RECT 0 86.975 0.070 88.725 ;
    RECT 0 88.795 0.070 90.545 ;
    RECT 0 90.615 0.070 92.365 ;
    RECT 0 92.435 0.070 94.185 ;
    RECT 0 94.255 0.070 96.005 ;
    RECT 0 96.075 0.070 97.825 ;
    RECT 0 97.895 0.070 99.645 ;
    RECT 0 99.715 0.070 101.465 ;
    RECT 0 101.535 0.070 103.285 ;
    RECT 0 103.355 0.070 105.105 ;
    RECT 0 105.175 0.070 106.925 ;
    RECT 0 106.995 0.070 108.745 ;
    RECT 0 108.815 0.070 110.565 ;
    RECT 0 110.635 0.070 112.385 ;
    RECT 0 112.455 0.070 114.205 ;
    RECT 0 114.275 0.070 116.025 ;
    RECT 0 116.095 0.070 117.845 ;
    RECT 0 117.915 0.070 119.665 ;
    RECT 0 119.735 0.070 121.485 ;
    RECT 0 121.555 0.070 123.305 ;
    RECT 0 123.375 0.070 125.125 ;
    RECT 0 125.195 0.070 126.945 ;
    RECT 0 127.015 0.070 128.765 ;
    RECT 0 128.835 0.070 130.585 ;
    RECT 0 130.655 0.070 132.405 ;
    RECT 0 132.475 0.070 134.225 ;
    RECT 0 134.295 0.070 136.045 ;
    RECT 0 136.115 0.070 137.865 ;
    RECT 0 137.935 0.070 139.685 ;
    RECT 0 139.755 0.070 141.505 ;
    RECT 0 141.575 0.070 143.325 ;
    RECT 0 143.395 0.070 145.145 ;
    RECT 0 145.215 0.070 146.965 ;
    RECT 0 147.035 0.070 148.785 ;
    RECT 0 148.855 0.070 150.605 ;
    RECT 0 150.675 0.070 152.425 ;
    RECT 0 152.495 0.070 154.245 ;
    RECT 0 154.315 0.070 156.065 ;
    RECT 0 156.135 0.070 157.885 ;
    RECT 0 157.955 0.070 159.705 ;
    RECT 0 159.775 0.070 161.525 ;
    RECT 0 161.595 0.070 163.345 ;
    RECT 0 163.415 0.070 165.165 ;
    RECT 0 165.235 0.070 166.985 ;
    RECT 0 167.055 0.070 168.805 ;
    RECT 0 168.875 0.070 170.625 ;
    RECT 0 170.695 0.070 172.445 ;
    RECT 0 172.515 0.070 174.265 ;
    RECT 0 174.335 0.070 178.745 ;
    RECT 0 178.815 0.070 180.565 ;
    RECT 0 180.635 0.070 182.385 ;
    RECT 0 182.455 0.070 184.205 ;
    RECT 0 184.275 0.070 186.025 ;
    RECT 0 186.095 0.070 187.845 ;
    RECT 0 187.915 0.070 189.665 ;
    RECT 0 189.735 0.070 191.485 ;
    RECT 0 191.555 0.070 193.305 ;
    RECT 0 193.375 0.070 195.125 ;
    RECT 0 195.195 0.070 196.945 ;
    RECT 0 197.015 0.070 198.765 ;
    RECT 0 198.835 0.070 200.585 ;
    RECT 0 200.655 0.070 202.405 ;
    RECT 0 202.475 0.070 204.225 ;
    RECT 0 204.295 0.070 206.045 ;
    RECT 0 206.115 0.070 207.865 ;
    RECT 0 207.935 0.070 209.685 ;
    RECT 0 209.755 0.070 211.505 ;
    RECT 0 211.575 0.070 213.325 ;
    RECT 0 213.395 0.070 215.145 ;
    RECT 0 215.215 0.070 216.965 ;
    RECT 0 217.035 0.070 218.785 ;
    RECT 0 218.855 0.070 220.605 ;
    RECT 0 220.675 0.070 222.425 ;
    RECT 0 222.495 0.070 224.245 ;
    RECT 0 224.315 0.070 226.065 ;
    RECT 0 226.135 0.070 227.885 ;
    RECT 0 227.955 0.070 229.705 ;
    RECT 0 229.775 0.070 231.525 ;
    RECT 0 231.595 0.070 233.345 ;
    RECT 0 233.415 0.070 235.165 ;
    RECT 0 235.235 0.070 236.985 ;
    RECT 0 237.055 0.070 238.805 ;
    RECT 0 238.875 0.070 240.625 ;
    RECT 0 240.695 0.070 242.445 ;
    RECT 0 242.515 0.070 244.265 ;
    RECT 0 244.335 0.070 246.085 ;
    RECT 0 246.155 0.070 247.905 ;
    RECT 0 247.975 0.070 249.725 ;
    RECT 0 249.795 0.070 251.545 ;
    RECT 0 251.615 0.070 253.365 ;
    RECT 0 253.435 0.070 255.185 ;
    RECT 0 255.255 0.070 257.005 ;
    RECT 0 257.075 0.070 258.825 ;
    RECT 0 258.895 0.070 260.645 ;
    RECT 0 260.715 0.070 262.465 ;
    RECT 0 262.535 0.070 264.285 ;
    RECT 0 264.355 0.070 266.105 ;
    RECT 0 266.175 0.070 267.925 ;
    RECT 0 267.995 0.070 269.745 ;
    RECT 0 269.815 0.070 271.565 ;
    RECT 0 271.635 0.070 273.385 ;
    RECT 0 273.455 0.070 275.205 ;
    RECT 0 275.275 0.070 277.025 ;
    RECT 0 277.095 0.070 278.845 ;
    RECT 0 278.915 0.070 280.665 ;
    RECT 0 280.735 0.070 282.485 ;
    RECT 0 282.555 0.070 284.305 ;
    RECT 0 284.375 0.070 286.125 ;
    RECT 0 286.195 0.070 287.945 ;
    RECT 0 288.015 0.070 289.765 ;
    RECT 0 289.835 0.070 291.585 ;
    RECT 0 291.655 0.070 293.405 ;
    RECT 0 293.475 0.070 295.225 ;
    RECT 0 295.295 0.070 297.045 ;
    RECT 0 297.115 0.070 298.865 ;
    RECT 0 298.935 0.070 300.685 ;
    RECT 0 300.755 0.070 302.505 ;
    RECT 0 302.575 0.070 304.325 ;
    RECT 0 304.395 0.070 306.145 ;
    RECT 0 306.215 0.070 307.965 ;
    RECT 0 308.035 0.070 309.785 ;
    RECT 0 309.855 0.070 311.605 ;
    RECT 0 311.675 0.070 313.425 ;
    RECT 0 313.495 0.070 315.245 ;
    RECT 0 315.315 0.070 317.065 ;
    RECT 0 317.135 0.070 318.885 ;
    RECT 0 318.955 0.070 320.705 ;
    RECT 0 320.775 0.070 322.525 ;
    RECT 0 322.595 0.070 324.345 ;
    RECT 0 324.415 0.070 326.165 ;
    RECT 0 326.235 0.070 327.985 ;
    RECT 0 328.055 0.070 329.805 ;
    RECT 0 329.875 0.070 331.625 ;
    RECT 0 331.695 0.070 333.445 ;
    RECT 0 333.515 0.070 335.265 ;
    RECT 0 335.335 0.070 337.085 ;
    RECT 0 337.155 0.070 338.905 ;
    RECT 0 338.975 0.070 340.725 ;
    RECT 0 340.795 0.070 342.545 ;
    RECT 0 342.615 0.070 344.365 ;
    RECT 0 344.435 0.070 346.185 ;
    RECT 0 346.255 0.070 348.005 ;
    RECT 0 348.075 0.070 349.825 ;
    RECT 0 349.895 0.070 351.645 ;
    RECT 0 351.715 0.070 356.125 ;
    RECT 0 356.195 0.070 357.945 ;
    RECT 0 358.015 0.070 359.765 ;
    RECT 0 359.835 0.070 361.585 ;
    RECT 0 361.655 0.070 363.405 ;
    RECT 0 363.475 0.070 365.225 ;
    RECT 0 365.295 0.070 367.045 ;
    RECT 0 367.115 0.070 368.865 ;
    RECT 0 368.935 0.070 370.685 ;
    RECT 0 370.755 0.070 372.505 ;
    RECT 0 372.575 0.070 374.325 ;
    RECT 0 374.395 0.070 376.145 ;
    RECT 0 376.215 0.070 377.965 ;
    RECT 0 378.035 0.070 379.785 ;
    RECT 0 379.855 0.070 381.605 ;
    RECT 0 381.675 0.070 383.425 ;
    RECT 0 383.495 0.070 385.245 ;
    RECT 0 385.315 0.070 387.065 ;
    RECT 0 387.135 0.070 388.885 ;
    RECT 0 388.955 0.070 390.705 ;
    RECT 0 390.775 0.070 392.525 ;
    RECT 0 392.595 0.070 394.345 ;
    RECT 0 394.415 0.070 396.165 ;
    RECT 0 396.235 0.070 397.985 ;
    RECT 0 398.055 0.070 399.805 ;
    RECT 0 399.875 0.070 401.625 ;
    RECT 0 401.695 0.070 403.445 ;
    RECT 0 403.515 0.070 405.265 ;
    RECT 0 405.335 0.070 407.085 ;
    RECT 0 407.155 0.070 408.905 ;
    RECT 0 408.975 0.070 410.725 ;
    RECT 0 410.795 0.070 412.545 ;
    RECT 0 412.615 0.070 414.365 ;
    RECT 0 414.435 0.070 416.185 ;
    RECT 0 416.255 0.070 418.005 ;
    RECT 0 418.075 0.070 419.825 ;
    RECT 0 419.895 0.070 421.645 ;
    RECT 0 421.715 0.070 423.465 ;
    RECT 0 423.535 0.070 425.285 ;
    RECT 0 425.355 0.070 427.105 ;
    RECT 0 427.175 0.070 428.925 ;
    RECT 0 428.995 0.070 430.745 ;
    RECT 0 430.815 0.070 432.565 ;
    RECT 0 432.635 0.070 434.385 ;
    RECT 0 434.455 0.070 436.205 ;
    RECT 0 436.275 0.070 438.025 ;
    RECT 0 438.095 0.070 439.845 ;
    RECT 0 439.915 0.070 441.665 ;
    RECT 0 441.735 0.070 443.485 ;
    RECT 0 443.555 0.070 445.305 ;
    RECT 0 445.375 0.070 447.125 ;
    RECT 0 447.195 0.070 448.945 ;
    RECT 0 449.015 0.070 450.765 ;
    RECT 0 450.835 0.070 452.585 ;
    RECT 0 452.655 0.070 454.405 ;
    RECT 0 454.475 0.070 456.225 ;
    RECT 0 456.295 0.070 458.045 ;
    RECT 0 458.115 0.070 459.865 ;
    RECT 0 459.935 0.070 461.685 ;
    RECT 0 461.755 0.070 463.505 ;
    RECT 0 463.575 0.070 465.325 ;
    RECT 0 465.395 0.070 467.145 ;
    RECT 0 467.215 0.070 468.965 ;
    RECT 0 469.035 0.070 470.785 ;
    RECT 0 470.855 0.070 472.605 ;
    RECT 0 472.675 0.070 474.425 ;
    RECT 0 474.495 0.070 476.245 ;
    RECT 0 476.315 0.070 478.065 ;
    RECT 0 478.135 0.070 479.885 ;
    RECT 0 479.955 0.070 481.705 ;
    RECT 0 481.775 0.070 483.525 ;
    RECT 0 483.595 0.070 485.345 ;
    RECT 0 485.415 0.070 487.165 ;
    RECT 0 487.235 0.070 488.985 ;
    RECT 0 489.055 0.070 490.805 ;
    RECT 0 490.875 0.070 492.625 ;
    RECT 0 492.695 0.070 494.445 ;
    RECT 0 494.515 0.070 496.265 ;
    RECT 0 496.335 0.070 498.085 ;
    RECT 0 498.155 0.070 499.905 ;
    RECT 0 499.975 0.070 501.725 ;
    RECT 0 501.795 0.070 503.545 ;
    RECT 0 503.615 0.070 505.365 ;
    RECT 0 505.435 0.070 507.185 ;
    RECT 0 507.255 0.070 509.005 ;
    RECT 0 509.075 0.070 510.825 ;
    RECT 0 510.895 0.070 512.645 ;
    RECT 0 512.715 0.070 514.465 ;
    RECT 0 514.535 0.070 516.285 ;
    RECT 0 516.355 0.070 518.105 ;
    RECT 0 518.175 0.070 519.925 ;
    RECT 0 519.995 0.070 521.745 ;
    RECT 0 521.815 0.070 523.565 ;
    RECT 0 523.635 0.070 525.385 ;
    RECT 0 525.455 0.070 527.205 ;
    RECT 0 527.275 0.070 529.025 ;
    RECT 0 529.095 0.070 533.505 ;
    RECT 0 533.575 0.070 535.325 ;
    RECT 0 535.395 0.070 537.145 ;
    RECT 0 537.215 0.070 538.965 ;
    RECT 0 539.035 0.070 540.785 ;
    RECT 0 540.855 0.070 542.605 ;
    RECT 0 542.675 0.070 544.425 ;
    RECT 0 544.495 0.070 546.245 ;
    RECT 0 546.315 0.070 548.065 ;
    RECT 0 548.135 0.070 549.885 ;
    RECT 0 549.955 0.070 551.705 ;
    RECT 0 551.775 0.070 553.525 ;
    RECT 0 553.595 0.070 558.005 ;
    RECT 0 558.075 0.070 559.825 ;
    RECT 0 559.895 0.070 561.645 ;
    RECT 0 561.715 0.070 572.600 ;
    LAYER metal4 ;
    RECT 0 0 747.080 1.400 ;
    RECT 0 571.200 747.080 572.600 ;
    RECT 0.000 1.400 1.260 571.200 ;
    RECT 1.540 1.400 2.380 571.200 ;
    RECT 2.660 1.400 3.500 571.200 ;
    RECT 3.780 1.400 4.620 571.200 ;
    RECT 4.900 1.400 5.740 571.200 ;
    RECT 6.020 1.400 6.860 571.200 ;
    RECT 7.140 1.400 7.980 571.200 ;
    RECT 8.260 1.400 9.100 571.200 ;
    RECT 9.380 1.400 10.220 571.200 ;
    RECT 10.500 1.400 11.340 571.200 ;
    RECT 11.620 1.400 12.460 571.200 ;
    RECT 12.740 1.400 13.580 571.200 ;
    RECT 13.860 1.400 14.700 571.200 ;
    RECT 14.980 1.400 15.820 571.200 ;
    RECT 16.100 1.400 16.940 571.200 ;
    RECT 17.220 1.400 18.060 571.200 ;
    RECT 18.340 1.400 19.180 571.200 ;
    RECT 19.460 1.400 20.300 571.200 ;
    RECT 20.580 1.400 21.420 571.200 ;
    RECT 21.700 1.400 22.540 571.200 ;
    RECT 22.820 1.400 23.660 571.200 ;
    RECT 23.940 1.400 24.780 571.200 ;
    RECT 25.060 1.400 25.900 571.200 ;
    RECT 26.180 1.400 27.020 571.200 ;
    RECT 27.300 1.400 28.140 571.200 ;
    RECT 28.420 1.400 29.260 571.200 ;
    RECT 29.540 1.400 30.380 571.200 ;
    RECT 30.660 1.400 31.500 571.200 ;
    RECT 31.780 1.400 32.620 571.200 ;
    RECT 32.900 1.400 33.740 571.200 ;
    RECT 34.020 1.400 34.860 571.200 ;
    RECT 35.140 1.400 35.980 571.200 ;
    RECT 36.260 1.400 37.100 571.200 ;
    RECT 37.380 1.400 38.220 571.200 ;
    RECT 38.500 1.400 39.340 571.200 ;
    RECT 39.620 1.400 40.460 571.200 ;
    RECT 40.740 1.400 41.580 571.200 ;
    RECT 41.860 1.400 42.700 571.200 ;
    RECT 42.980 1.400 43.820 571.200 ;
    RECT 44.100 1.400 44.940 571.200 ;
    RECT 45.220 1.400 46.060 571.200 ;
    RECT 46.340 1.400 47.180 571.200 ;
    RECT 47.460 1.400 48.300 571.200 ;
    RECT 48.580 1.400 49.420 571.200 ;
    RECT 49.700 1.400 50.540 571.200 ;
    RECT 50.820 1.400 51.660 571.200 ;
    RECT 51.940 1.400 52.780 571.200 ;
    RECT 53.060 1.400 53.900 571.200 ;
    RECT 54.180 1.400 55.020 571.200 ;
    RECT 55.300 1.400 56.140 571.200 ;
    RECT 56.420 1.400 57.260 571.200 ;
    RECT 57.540 1.400 58.380 571.200 ;
    RECT 58.660 1.400 59.500 571.200 ;
    RECT 59.780 1.400 60.620 571.200 ;
    RECT 60.900 1.400 61.740 571.200 ;
    RECT 62.020 1.400 62.860 571.200 ;
    RECT 63.140 1.400 63.980 571.200 ;
    RECT 64.260 1.400 65.100 571.200 ;
    RECT 65.380 1.400 66.220 571.200 ;
    RECT 66.500 1.400 67.340 571.200 ;
    RECT 67.620 1.400 68.460 571.200 ;
    RECT 68.740 1.400 69.580 571.200 ;
    RECT 69.860 1.400 70.700 571.200 ;
    RECT 70.980 1.400 71.820 571.200 ;
    RECT 72.100 1.400 72.940 571.200 ;
    RECT 73.220 1.400 74.060 571.200 ;
    RECT 74.340 1.400 75.180 571.200 ;
    RECT 75.460 1.400 76.300 571.200 ;
    RECT 76.580 1.400 77.420 571.200 ;
    RECT 77.700 1.400 78.540 571.200 ;
    RECT 78.820 1.400 79.660 571.200 ;
    RECT 79.940 1.400 80.780 571.200 ;
    RECT 81.060 1.400 81.900 571.200 ;
    RECT 82.180 1.400 83.020 571.200 ;
    RECT 83.300 1.400 84.140 571.200 ;
    RECT 84.420 1.400 85.260 571.200 ;
    RECT 85.540 1.400 86.380 571.200 ;
    RECT 86.660 1.400 87.500 571.200 ;
    RECT 87.780 1.400 88.620 571.200 ;
    RECT 88.900 1.400 89.740 571.200 ;
    RECT 90.020 1.400 90.860 571.200 ;
    RECT 91.140 1.400 91.980 571.200 ;
    RECT 92.260 1.400 93.100 571.200 ;
    RECT 93.380 1.400 94.220 571.200 ;
    RECT 94.500 1.400 95.340 571.200 ;
    RECT 95.620 1.400 96.460 571.200 ;
    RECT 96.740 1.400 97.580 571.200 ;
    RECT 97.860 1.400 98.700 571.200 ;
    RECT 98.980 1.400 99.820 571.200 ;
    RECT 100.100 1.400 100.940 571.200 ;
    RECT 101.220 1.400 102.060 571.200 ;
    RECT 102.340 1.400 103.180 571.200 ;
    RECT 103.460 1.400 104.300 571.200 ;
    RECT 104.580 1.400 105.420 571.200 ;
    RECT 105.700 1.400 106.540 571.200 ;
    RECT 106.820 1.400 107.660 571.200 ;
    RECT 107.940 1.400 108.780 571.200 ;
    RECT 109.060 1.400 109.900 571.200 ;
    RECT 110.180 1.400 111.020 571.200 ;
    RECT 111.300 1.400 112.140 571.200 ;
    RECT 112.420 1.400 113.260 571.200 ;
    RECT 113.540 1.400 114.380 571.200 ;
    RECT 114.660 1.400 115.500 571.200 ;
    RECT 115.780 1.400 116.620 571.200 ;
    RECT 116.900 1.400 117.740 571.200 ;
    RECT 118.020 1.400 118.860 571.200 ;
    RECT 119.140 1.400 119.980 571.200 ;
    RECT 120.260 1.400 121.100 571.200 ;
    RECT 121.380 1.400 122.220 571.200 ;
    RECT 122.500 1.400 123.340 571.200 ;
    RECT 123.620 1.400 124.460 571.200 ;
    RECT 124.740 1.400 125.580 571.200 ;
    RECT 125.860 1.400 126.700 571.200 ;
    RECT 126.980 1.400 127.820 571.200 ;
    RECT 128.100 1.400 128.940 571.200 ;
    RECT 129.220 1.400 130.060 571.200 ;
    RECT 130.340 1.400 131.180 571.200 ;
    RECT 131.460 1.400 132.300 571.200 ;
    RECT 132.580 1.400 133.420 571.200 ;
    RECT 133.700 1.400 134.540 571.200 ;
    RECT 134.820 1.400 135.660 571.200 ;
    RECT 135.940 1.400 136.780 571.200 ;
    RECT 137.060 1.400 137.900 571.200 ;
    RECT 138.180 1.400 139.020 571.200 ;
    RECT 139.300 1.400 140.140 571.200 ;
    RECT 140.420 1.400 141.260 571.200 ;
    RECT 141.540 1.400 142.380 571.200 ;
    RECT 142.660 1.400 143.500 571.200 ;
    RECT 143.780 1.400 144.620 571.200 ;
    RECT 144.900 1.400 145.740 571.200 ;
    RECT 146.020 1.400 146.860 571.200 ;
    RECT 147.140 1.400 147.980 571.200 ;
    RECT 148.260 1.400 149.100 571.200 ;
    RECT 149.380 1.400 150.220 571.200 ;
    RECT 150.500 1.400 151.340 571.200 ;
    RECT 151.620 1.400 152.460 571.200 ;
    RECT 152.740 1.400 153.580 571.200 ;
    RECT 153.860 1.400 154.700 571.200 ;
    RECT 154.980 1.400 155.820 571.200 ;
    RECT 156.100 1.400 156.940 571.200 ;
    RECT 157.220 1.400 158.060 571.200 ;
    RECT 158.340 1.400 159.180 571.200 ;
    RECT 159.460 1.400 160.300 571.200 ;
    RECT 160.580 1.400 161.420 571.200 ;
    RECT 161.700 1.400 162.540 571.200 ;
    RECT 162.820 1.400 163.660 571.200 ;
    RECT 163.940 1.400 164.780 571.200 ;
    RECT 165.060 1.400 165.900 571.200 ;
    RECT 166.180 1.400 167.020 571.200 ;
    RECT 167.300 1.400 168.140 571.200 ;
    RECT 168.420 1.400 169.260 571.200 ;
    RECT 169.540 1.400 170.380 571.200 ;
    RECT 170.660 1.400 171.500 571.200 ;
    RECT 171.780 1.400 172.620 571.200 ;
    RECT 172.900 1.400 173.740 571.200 ;
    RECT 174.020 1.400 174.860 571.200 ;
    RECT 175.140 1.400 175.980 571.200 ;
    RECT 176.260 1.400 177.100 571.200 ;
    RECT 177.380 1.400 178.220 571.200 ;
    RECT 178.500 1.400 179.340 571.200 ;
    RECT 179.620 1.400 180.460 571.200 ;
    RECT 180.740 1.400 181.580 571.200 ;
    RECT 181.860 1.400 182.700 571.200 ;
    RECT 182.980 1.400 183.820 571.200 ;
    RECT 184.100 1.400 184.940 571.200 ;
    RECT 185.220 1.400 186.060 571.200 ;
    RECT 186.340 1.400 187.180 571.200 ;
    RECT 187.460 1.400 188.300 571.200 ;
    RECT 188.580 1.400 189.420 571.200 ;
    RECT 189.700 1.400 190.540 571.200 ;
    RECT 190.820 1.400 191.660 571.200 ;
    RECT 191.940 1.400 192.780 571.200 ;
    RECT 193.060 1.400 193.900 571.200 ;
    RECT 194.180 1.400 195.020 571.200 ;
    RECT 195.300 1.400 196.140 571.200 ;
    RECT 196.420 1.400 197.260 571.200 ;
    RECT 197.540 1.400 198.380 571.200 ;
    RECT 198.660 1.400 199.500 571.200 ;
    RECT 199.780 1.400 200.620 571.200 ;
    RECT 200.900 1.400 201.740 571.200 ;
    RECT 202.020 1.400 202.860 571.200 ;
    RECT 203.140 1.400 203.980 571.200 ;
    RECT 204.260 1.400 205.100 571.200 ;
    RECT 205.380 1.400 206.220 571.200 ;
    RECT 206.500 1.400 207.340 571.200 ;
    RECT 207.620 1.400 208.460 571.200 ;
    RECT 208.740 1.400 209.580 571.200 ;
    RECT 209.860 1.400 210.700 571.200 ;
    RECT 210.980 1.400 211.820 571.200 ;
    RECT 212.100 1.400 212.940 571.200 ;
    RECT 213.220 1.400 214.060 571.200 ;
    RECT 214.340 1.400 215.180 571.200 ;
    RECT 215.460 1.400 216.300 571.200 ;
    RECT 216.580 1.400 217.420 571.200 ;
    RECT 217.700 1.400 218.540 571.200 ;
    RECT 218.820 1.400 219.660 571.200 ;
    RECT 219.940 1.400 220.780 571.200 ;
    RECT 221.060 1.400 221.900 571.200 ;
    RECT 222.180 1.400 223.020 571.200 ;
    RECT 223.300 1.400 224.140 571.200 ;
    RECT 224.420 1.400 225.260 571.200 ;
    RECT 225.540 1.400 226.380 571.200 ;
    RECT 226.660 1.400 227.500 571.200 ;
    RECT 227.780 1.400 228.620 571.200 ;
    RECT 228.900 1.400 229.740 571.200 ;
    RECT 230.020 1.400 230.860 571.200 ;
    RECT 231.140 1.400 231.980 571.200 ;
    RECT 232.260 1.400 233.100 571.200 ;
    RECT 233.380 1.400 234.220 571.200 ;
    RECT 234.500 1.400 235.340 571.200 ;
    RECT 235.620 1.400 236.460 571.200 ;
    RECT 236.740 1.400 237.580 571.200 ;
    RECT 237.860 1.400 238.700 571.200 ;
    RECT 238.980 1.400 239.820 571.200 ;
    RECT 240.100 1.400 240.940 571.200 ;
    RECT 241.220 1.400 242.060 571.200 ;
    RECT 242.340 1.400 243.180 571.200 ;
    RECT 243.460 1.400 244.300 571.200 ;
    RECT 244.580 1.400 245.420 571.200 ;
    RECT 245.700 1.400 246.540 571.200 ;
    RECT 246.820 1.400 247.660 571.200 ;
    RECT 247.940 1.400 248.780 571.200 ;
    RECT 249.060 1.400 249.900 571.200 ;
    RECT 250.180 1.400 251.020 571.200 ;
    RECT 251.300 1.400 252.140 571.200 ;
    RECT 252.420 1.400 253.260 571.200 ;
    RECT 253.540 1.400 254.380 571.200 ;
    RECT 254.660 1.400 255.500 571.200 ;
    RECT 255.780 1.400 256.620 571.200 ;
    RECT 256.900 1.400 257.740 571.200 ;
    RECT 258.020 1.400 258.860 571.200 ;
    RECT 259.140 1.400 259.980 571.200 ;
    RECT 260.260 1.400 261.100 571.200 ;
    RECT 261.380 1.400 262.220 571.200 ;
    RECT 262.500 1.400 263.340 571.200 ;
    RECT 263.620 1.400 264.460 571.200 ;
    RECT 264.740 1.400 265.580 571.200 ;
    RECT 265.860 1.400 266.700 571.200 ;
    RECT 266.980 1.400 267.820 571.200 ;
    RECT 268.100 1.400 268.940 571.200 ;
    RECT 269.220 1.400 270.060 571.200 ;
    RECT 270.340 1.400 271.180 571.200 ;
    RECT 271.460 1.400 272.300 571.200 ;
    RECT 272.580 1.400 273.420 571.200 ;
    RECT 273.700 1.400 274.540 571.200 ;
    RECT 274.820 1.400 275.660 571.200 ;
    RECT 275.940 1.400 276.780 571.200 ;
    RECT 277.060 1.400 277.900 571.200 ;
    RECT 278.180 1.400 279.020 571.200 ;
    RECT 279.300 1.400 280.140 571.200 ;
    RECT 280.420 1.400 281.260 571.200 ;
    RECT 281.540 1.400 282.380 571.200 ;
    RECT 282.660 1.400 283.500 571.200 ;
    RECT 283.780 1.400 284.620 571.200 ;
    RECT 284.900 1.400 285.740 571.200 ;
    RECT 286.020 1.400 286.860 571.200 ;
    RECT 287.140 1.400 287.980 571.200 ;
    RECT 288.260 1.400 289.100 571.200 ;
    RECT 289.380 1.400 290.220 571.200 ;
    RECT 290.500 1.400 291.340 571.200 ;
    RECT 291.620 1.400 292.460 571.200 ;
    RECT 292.740 1.400 293.580 571.200 ;
    RECT 293.860 1.400 294.700 571.200 ;
    RECT 294.980 1.400 295.820 571.200 ;
    RECT 296.100 1.400 296.940 571.200 ;
    RECT 297.220 1.400 298.060 571.200 ;
    RECT 298.340 1.400 299.180 571.200 ;
    RECT 299.460 1.400 300.300 571.200 ;
    RECT 300.580 1.400 301.420 571.200 ;
    RECT 301.700 1.400 302.540 571.200 ;
    RECT 302.820 1.400 303.660 571.200 ;
    RECT 303.940 1.400 304.780 571.200 ;
    RECT 305.060 1.400 305.900 571.200 ;
    RECT 306.180 1.400 307.020 571.200 ;
    RECT 307.300 1.400 308.140 571.200 ;
    RECT 308.420 1.400 309.260 571.200 ;
    RECT 309.540 1.400 310.380 571.200 ;
    RECT 310.660 1.400 311.500 571.200 ;
    RECT 311.780 1.400 312.620 571.200 ;
    RECT 312.900 1.400 313.740 571.200 ;
    RECT 314.020 1.400 314.860 571.200 ;
    RECT 315.140 1.400 315.980 571.200 ;
    RECT 316.260 1.400 317.100 571.200 ;
    RECT 317.380 1.400 318.220 571.200 ;
    RECT 318.500 1.400 319.340 571.200 ;
    RECT 319.620 1.400 320.460 571.200 ;
    RECT 320.740 1.400 321.580 571.200 ;
    RECT 321.860 1.400 322.700 571.200 ;
    RECT 322.980 1.400 323.820 571.200 ;
    RECT 324.100 1.400 324.940 571.200 ;
    RECT 325.220 1.400 326.060 571.200 ;
    RECT 326.340 1.400 327.180 571.200 ;
    RECT 327.460 1.400 328.300 571.200 ;
    RECT 328.580 1.400 329.420 571.200 ;
    RECT 329.700 1.400 330.540 571.200 ;
    RECT 330.820 1.400 331.660 571.200 ;
    RECT 331.940 1.400 332.780 571.200 ;
    RECT 333.060 1.400 333.900 571.200 ;
    RECT 334.180 1.400 335.020 571.200 ;
    RECT 335.300 1.400 336.140 571.200 ;
    RECT 336.420 1.400 337.260 571.200 ;
    RECT 337.540 1.400 338.380 571.200 ;
    RECT 338.660 1.400 339.500 571.200 ;
    RECT 339.780 1.400 340.620 571.200 ;
    RECT 340.900 1.400 341.740 571.200 ;
    RECT 342.020 1.400 342.860 571.200 ;
    RECT 343.140 1.400 343.980 571.200 ;
    RECT 344.260 1.400 345.100 571.200 ;
    RECT 345.380 1.400 346.220 571.200 ;
    RECT 346.500 1.400 347.340 571.200 ;
    RECT 347.620 1.400 348.460 571.200 ;
    RECT 348.740 1.400 349.580 571.200 ;
    RECT 349.860 1.400 350.700 571.200 ;
    RECT 350.980 1.400 351.820 571.200 ;
    RECT 352.100 1.400 352.940 571.200 ;
    RECT 353.220 1.400 354.060 571.200 ;
    RECT 354.340 1.400 355.180 571.200 ;
    RECT 355.460 1.400 356.300 571.200 ;
    RECT 356.580 1.400 357.420 571.200 ;
    RECT 357.700 1.400 358.540 571.200 ;
    RECT 358.820 1.400 359.660 571.200 ;
    RECT 359.940 1.400 360.780 571.200 ;
    RECT 361.060 1.400 361.900 571.200 ;
    RECT 362.180 1.400 363.020 571.200 ;
    RECT 363.300 1.400 364.140 571.200 ;
    RECT 364.420 1.400 365.260 571.200 ;
    RECT 365.540 1.400 366.380 571.200 ;
    RECT 366.660 1.400 367.500 571.200 ;
    RECT 367.780 1.400 368.620 571.200 ;
    RECT 368.900 1.400 369.740 571.200 ;
    RECT 370.020 1.400 370.860 571.200 ;
    RECT 371.140 1.400 371.980 571.200 ;
    RECT 372.260 1.400 373.100 571.200 ;
    RECT 373.380 1.400 374.220 571.200 ;
    RECT 374.500 1.400 375.340 571.200 ;
    RECT 375.620 1.400 376.460 571.200 ;
    RECT 376.740 1.400 377.580 571.200 ;
    RECT 377.860 1.400 378.700 571.200 ;
    RECT 378.980 1.400 379.820 571.200 ;
    RECT 380.100 1.400 380.940 571.200 ;
    RECT 381.220 1.400 382.060 571.200 ;
    RECT 382.340 1.400 383.180 571.200 ;
    RECT 383.460 1.400 384.300 571.200 ;
    RECT 384.580 1.400 385.420 571.200 ;
    RECT 385.700 1.400 386.540 571.200 ;
    RECT 386.820 1.400 387.660 571.200 ;
    RECT 387.940 1.400 388.780 571.200 ;
    RECT 389.060 1.400 389.900 571.200 ;
    RECT 390.180 1.400 391.020 571.200 ;
    RECT 391.300 1.400 392.140 571.200 ;
    RECT 392.420 1.400 393.260 571.200 ;
    RECT 393.540 1.400 394.380 571.200 ;
    RECT 394.660 1.400 395.500 571.200 ;
    RECT 395.780 1.400 396.620 571.200 ;
    RECT 396.900 1.400 397.740 571.200 ;
    RECT 398.020 1.400 398.860 571.200 ;
    RECT 399.140 1.400 399.980 571.200 ;
    RECT 400.260 1.400 401.100 571.200 ;
    RECT 401.380 1.400 402.220 571.200 ;
    RECT 402.500 1.400 403.340 571.200 ;
    RECT 403.620 1.400 404.460 571.200 ;
    RECT 404.740 1.400 405.580 571.200 ;
    RECT 405.860 1.400 406.700 571.200 ;
    RECT 406.980 1.400 407.820 571.200 ;
    RECT 408.100 1.400 408.940 571.200 ;
    RECT 409.220 1.400 410.060 571.200 ;
    RECT 410.340 1.400 411.180 571.200 ;
    RECT 411.460 1.400 412.300 571.200 ;
    RECT 412.580 1.400 413.420 571.200 ;
    RECT 413.700 1.400 414.540 571.200 ;
    RECT 414.820 1.400 415.660 571.200 ;
    RECT 415.940 1.400 416.780 571.200 ;
    RECT 417.060 1.400 417.900 571.200 ;
    RECT 418.180 1.400 419.020 571.200 ;
    RECT 419.300 1.400 420.140 571.200 ;
    RECT 420.420 1.400 421.260 571.200 ;
    RECT 421.540 1.400 422.380 571.200 ;
    RECT 422.660 1.400 423.500 571.200 ;
    RECT 423.780 1.400 424.620 571.200 ;
    RECT 424.900 1.400 425.740 571.200 ;
    RECT 426.020 1.400 426.860 571.200 ;
    RECT 427.140 1.400 427.980 571.200 ;
    RECT 428.260 1.400 429.100 571.200 ;
    RECT 429.380 1.400 430.220 571.200 ;
    RECT 430.500 1.400 431.340 571.200 ;
    RECT 431.620 1.400 432.460 571.200 ;
    RECT 432.740 1.400 433.580 571.200 ;
    RECT 433.860 1.400 434.700 571.200 ;
    RECT 434.980 1.400 435.820 571.200 ;
    RECT 436.100 1.400 436.940 571.200 ;
    RECT 437.220 1.400 438.060 571.200 ;
    RECT 438.340 1.400 439.180 571.200 ;
    RECT 439.460 1.400 440.300 571.200 ;
    RECT 440.580 1.400 441.420 571.200 ;
    RECT 441.700 1.400 442.540 571.200 ;
    RECT 442.820 1.400 443.660 571.200 ;
    RECT 443.940 1.400 444.780 571.200 ;
    RECT 445.060 1.400 445.900 571.200 ;
    RECT 446.180 1.400 447.020 571.200 ;
    RECT 447.300 1.400 448.140 571.200 ;
    RECT 448.420 1.400 449.260 571.200 ;
    RECT 449.540 1.400 450.380 571.200 ;
    RECT 450.660 1.400 451.500 571.200 ;
    RECT 451.780 1.400 452.620 571.200 ;
    RECT 452.900 1.400 453.740 571.200 ;
    RECT 454.020 1.400 454.860 571.200 ;
    RECT 455.140 1.400 455.980 571.200 ;
    RECT 456.260 1.400 457.100 571.200 ;
    RECT 457.380 1.400 458.220 571.200 ;
    RECT 458.500 1.400 459.340 571.200 ;
    RECT 459.620 1.400 460.460 571.200 ;
    RECT 460.740 1.400 461.580 571.200 ;
    RECT 461.860 1.400 462.700 571.200 ;
    RECT 462.980 1.400 463.820 571.200 ;
    RECT 464.100 1.400 464.940 571.200 ;
    RECT 465.220 1.400 466.060 571.200 ;
    RECT 466.340 1.400 467.180 571.200 ;
    RECT 467.460 1.400 468.300 571.200 ;
    RECT 468.580 1.400 469.420 571.200 ;
    RECT 469.700 1.400 470.540 571.200 ;
    RECT 470.820 1.400 471.660 571.200 ;
    RECT 471.940 1.400 472.780 571.200 ;
    RECT 473.060 1.400 473.900 571.200 ;
    RECT 474.180 1.400 475.020 571.200 ;
    RECT 475.300 1.400 476.140 571.200 ;
    RECT 476.420 1.400 477.260 571.200 ;
    RECT 477.540 1.400 478.380 571.200 ;
    RECT 478.660 1.400 479.500 571.200 ;
    RECT 479.780 1.400 480.620 571.200 ;
    RECT 480.900 1.400 481.740 571.200 ;
    RECT 482.020 1.400 482.860 571.200 ;
    RECT 483.140 1.400 483.980 571.200 ;
    RECT 484.260 1.400 485.100 571.200 ;
    RECT 485.380 1.400 486.220 571.200 ;
    RECT 486.500 1.400 487.340 571.200 ;
    RECT 487.620 1.400 488.460 571.200 ;
    RECT 488.740 1.400 489.580 571.200 ;
    RECT 489.860 1.400 490.700 571.200 ;
    RECT 490.980 1.400 491.820 571.200 ;
    RECT 492.100 1.400 492.940 571.200 ;
    RECT 493.220 1.400 494.060 571.200 ;
    RECT 494.340 1.400 495.180 571.200 ;
    RECT 495.460 1.400 496.300 571.200 ;
    RECT 496.580 1.400 497.420 571.200 ;
    RECT 497.700 1.400 498.540 571.200 ;
    RECT 498.820 1.400 499.660 571.200 ;
    RECT 499.940 1.400 500.780 571.200 ;
    RECT 501.060 1.400 501.900 571.200 ;
    RECT 502.180 1.400 503.020 571.200 ;
    RECT 503.300 1.400 504.140 571.200 ;
    RECT 504.420 1.400 505.260 571.200 ;
    RECT 505.540 1.400 506.380 571.200 ;
    RECT 506.660 1.400 507.500 571.200 ;
    RECT 507.780 1.400 508.620 571.200 ;
    RECT 508.900 1.400 509.740 571.200 ;
    RECT 510.020 1.400 510.860 571.200 ;
    RECT 511.140 1.400 511.980 571.200 ;
    RECT 512.260 1.400 513.100 571.200 ;
    RECT 513.380 1.400 514.220 571.200 ;
    RECT 514.500 1.400 515.340 571.200 ;
    RECT 515.620 1.400 516.460 571.200 ;
    RECT 516.740 1.400 517.580 571.200 ;
    RECT 517.860 1.400 518.700 571.200 ;
    RECT 518.980 1.400 519.820 571.200 ;
    RECT 520.100 1.400 520.940 571.200 ;
    RECT 521.220 1.400 522.060 571.200 ;
    RECT 522.340 1.400 523.180 571.200 ;
    RECT 523.460 1.400 524.300 571.200 ;
    RECT 524.580 1.400 525.420 571.200 ;
    RECT 525.700 1.400 526.540 571.200 ;
    RECT 526.820 1.400 527.660 571.200 ;
    RECT 527.940 1.400 528.780 571.200 ;
    RECT 529.060 1.400 529.900 571.200 ;
    RECT 530.180 1.400 531.020 571.200 ;
    RECT 531.300 1.400 532.140 571.200 ;
    RECT 532.420 1.400 533.260 571.200 ;
    RECT 533.540 1.400 534.380 571.200 ;
    RECT 534.660 1.400 535.500 571.200 ;
    RECT 535.780 1.400 536.620 571.200 ;
    RECT 536.900 1.400 537.740 571.200 ;
    RECT 538.020 1.400 538.860 571.200 ;
    RECT 539.140 1.400 539.980 571.200 ;
    RECT 540.260 1.400 541.100 571.200 ;
    RECT 541.380 1.400 542.220 571.200 ;
    RECT 542.500 1.400 543.340 571.200 ;
    RECT 543.620 1.400 544.460 571.200 ;
    RECT 544.740 1.400 545.580 571.200 ;
    RECT 545.860 1.400 546.700 571.200 ;
    RECT 546.980 1.400 547.820 571.200 ;
    RECT 548.100 1.400 548.940 571.200 ;
    RECT 549.220 1.400 550.060 571.200 ;
    RECT 550.340 1.400 551.180 571.200 ;
    RECT 551.460 1.400 552.300 571.200 ;
    RECT 552.580 1.400 553.420 571.200 ;
    RECT 553.700 1.400 554.540 571.200 ;
    RECT 554.820 1.400 555.660 571.200 ;
    RECT 555.940 1.400 556.780 571.200 ;
    RECT 557.060 1.400 557.900 571.200 ;
    RECT 558.180 1.400 559.020 571.200 ;
    RECT 559.300 1.400 560.140 571.200 ;
    RECT 560.420 1.400 561.260 571.200 ;
    RECT 561.540 1.400 562.380 571.200 ;
    RECT 562.660 1.400 563.500 571.200 ;
    RECT 563.780 1.400 564.620 571.200 ;
    RECT 564.900 1.400 565.740 571.200 ;
    RECT 566.020 1.400 566.860 571.200 ;
    RECT 567.140 1.400 567.980 571.200 ;
    RECT 568.260 1.400 569.100 571.200 ;
    RECT 569.380 1.400 570.220 571.200 ;
    RECT 570.500 1.400 571.340 571.200 ;
    RECT 571.620 1.400 572.460 571.200 ;
    RECT 572.740 1.400 573.580 571.200 ;
    RECT 573.860 1.400 574.700 571.200 ;
    RECT 574.980 1.400 575.820 571.200 ;
    RECT 576.100 1.400 576.940 571.200 ;
    RECT 577.220 1.400 578.060 571.200 ;
    RECT 578.340 1.400 579.180 571.200 ;
    RECT 579.460 1.400 580.300 571.200 ;
    RECT 580.580 1.400 581.420 571.200 ;
    RECT 581.700 1.400 582.540 571.200 ;
    RECT 582.820 1.400 583.660 571.200 ;
    RECT 583.940 1.400 584.780 571.200 ;
    RECT 585.060 1.400 585.900 571.200 ;
    RECT 586.180 1.400 587.020 571.200 ;
    RECT 587.300 1.400 588.140 571.200 ;
    RECT 588.420 1.400 589.260 571.200 ;
    RECT 589.540 1.400 590.380 571.200 ;
    RECT 590.660 1.400 591.500 571.200 ;
    RECT 591.780 1.400 592.620 571.200 ;
    RECT 592.900 1.400 593.740 571.200 ;
    RECT 594.020 1.400 594.860 571.200 ;
    RECT 595.140 1.400 595.980 571.200 ;
    RECT 596.260 1.400 597.100 571.200 ;
    RECT 597.380 1.400 598.220 571.200 ;
    RECT 598.500 1.400 599.340 571.200 ;
    RECT 599.620 1.400 600.460 571.200 ;
    RECT 600.740 1.400 601.580 571.200 ;
    RECT 601.860 1.400 602.700 571.200 ;
    RECT 602.980 1.400 603.820 571.200 ;
    RECT 604.100 1.400 604.940 571.200 ;
    RECT 605.220 1.400 606.060 571.200 ;
    RECT 606.340 1.400 607.180 571.200 ;
    RECT 607.460 1.400 608.300 571.200 ;
    RECT 608.580 1.400 609.420 571.200 ;
    RECT 609.700 1.400 610.540 571.200 ;
    RECT 610.820 1.400 611.660 571.200 ;
    RECT 611.940 1.400 612.780 571.200 ;
    RECT 613.060 1.400 613.900 571.200 ;
    RECT 614.180 1.400 615.020 571.200 ;
    RECT 615.300 1.400 616.140 571.200 ;
    RECT 616.420 1.400 617.260 571.200 ;
    RECT 617.540 1.400 618.380 571.200 ;
    RECT 618.660 1.400 619.500 571.200 ;
    RECT 619.780 1.400 620.620 571.200 ;
    RECT 620.900 1.400 621.740 571.200 ;
    RECT 622.020 1.400 622.860 571.200 ;
    RECT 623.140 1.400 623.980 571.200 ;
    RECT 624.260 1.400 625.100 571.200 ;
    RECT 625.380 1.400 626.220 571.200 ;
    RECT 626.500 1.400 627.340 571.200 ;
    RECT 627.620 1.400 628.460 571.200 ;
    RECT 628.740 1.400 629.580 571.200 ;
    RECT 629.860 1.400 630.700 571.200 ;
    RECT 630.980 1.400 631.820 571.200 ;
    RECT 632.100 1.400 632.940 571.200 ;
    RECT 633.220 1.400 634.060 571.200 ;
    RECT 634.340 1.400 635.180 571.200 ;
    RECT 635.460 1.400 636.300 571.200 ;
    RECT 636.580 1.400 637.420 571.200 ;
    RECT 637.700 1.400 638.540 571.200 ;
    RECT 638.820 1.400 639.660 571.200 ;
    RECT 639.940 1.400 640.780 571.200 ;
    RECT 641.060 1.400 641.900 571.200 ;
    RECT 642.180 1.400 643.020 571.200 ;
    RECT 643.300 1.400 644.140 571.200 ;
    RECT 644.420 1.400 645.260 571.200 ;
    RECT 645.540 1.400 646.380 571.200 ;
    RECT 646.660 1.400 647.500 571.200 ;
    RECT 647.780 1.400 648.620 571.200 ;
    RECT 648.900 1.400 649.740 571.200 ;
    RECT 650.020 1.400 650.860 571.200 ;
    RECT 651.140 1.400 651.980 571.200 ;
    RECT 652.260 1.400 653.100 571.200 ;
    RECT 653.380 1.400 654.220 571.200 ;
    RECT 654.500 1.400 655.340 571.200 ;
    RECT 655.620 1.400 656.460 571.200 ;
    RECT 656.740 1.400 657.580 571.200 ;
    RECT 657.860 1.400 658.700 571.200 ;
    RECT 658.980 1.400 659.820 571.200 ;
    RECT 660.100 1.400 660.940 571.200 ;
    RECT 661.220 1.400 662.060 571.200 ;
    RECT 662.340 1.400 663.180 571.200 ;
    RECT 663.460 1.400 664.300 571.200 ;
    RECT 664.580 1.400 665.420 571.200 ;
    RECT 665.700 1.400 666.540 571.200 ;
    RECT 666.820 1.400 667.660 571.200 ;
    RECT 667.940 1.400 668.780 571.200 ;
    RECT 669.060 1.400 669.900 571.200 ;
    RECT 670.180 1.400 671.020 571.200 ;
    RECT 671.300 1.400 672.140 571.200 ;
    RECT 672.420 1.400 673.260 571.200 ;
    RECT 673.540 1.400 674.380 571.200 ;
    RECT 674.660 1.400 675.500 571.200 ;
    RECT 675.780 1.400 676.620 571.200 ;
    RECT 676.900 1.400 677.740 571.200 ;
    RECT 678.020 1.400 678.860 571.200 ;
    RECT 679.140 1.400 679.980 571.200 ;
    RECT 680.260 1.400 681.100 571.200 ;
    RECT 681.380 1.400 682.220 571.200 ;
    RECT 682.500 1.400 683.340 571.200 ;
    RECT 683.620 1.400 684.460 571.200 ;
    RECT 684.740 1.400 685.580 571.200 ;
    RECT 685.860 1.400 686.700 571.200 ;
    RECT 686.980 1.400 687.820 571.200 ;
    RECT 688.100 1.400 688.940 571.200 ;
    RECT 689.220 1.400 690.060 571.200 ;
    RECT 690.340 1.400 691.180 571.200 ;
    RECT 691.460 1.400 692.300 571.200 ;
    RECT 692.580 1.400 693.420 571.200 ;
    RECT 693.700 1.400 694.540 571.200 ;
    RECT 694.820 1.400 695.660 571.200 ;
    RECT 695.940 1.400 696.780 571.200 ;
    RECT 697.060 1.400 697.900 571.200 ;
    RECT 698.180 1.400 699.020 571.200 ;
    RECT 699.300 1.400 700.140 571.200 ;
    RECT 700.420 1.400 701.260 571.200 ;
    RECT 701.540 1.400 702.380 571.200 ;
    RECT 702.660 1.400 703.500 571.200 ;
    RECT 703.780 1.400 704.620 571.200 ;
    RECT 704.900 1.400 705.740 571.200 ;
    RECT 706.020 1.400 706.860 571.200 ;
    RECT 707.140 1.400 707.980 571.200 ;
    RECT 708.260 1.400 709.100 571.200 ;
    RECT 709.380 1.400 710.220 571.200 ;
    RECT 710.500 1.400 711.340 571.200 ;
    RECT 711.620 1.400 712.460 571.200 ;
    RECT 712.740 1.400 713.580 571.200 ;
    RECT 713.860 1.400 714.700 571.200 ;
    RECT 714.980 1.400 715.820 571.200 ;
    RECT 716.100 1.400 716.940 571.200 ;
    RECT 717.220 1.400 718.060 571.200 ;
    RECT 718.340 1.400 719.180 571.200 ;
    RECT 719.460 1.400 720.300 571.200 ;
    RECT 720.580 1.400 721.420 571.200 ;
    RECT 721.700 1.400 722.540 571.200 ;
    RECT 722.820 1.400 723.660 571.200 ;
    RECT 723.940 1.400 724.780 571.200 ;
    RECT 725.060 1.400 725.900 571.200 ;
    RECT 726.180 1.400 727.020 571.200 ;
    RECT 727.300 1.400 728.140 571.200 ;
    RECT 728.420 1.400 729.260 571.200 ;
    RECT 729.540 1.400 730.380 571.200 ;
    RECT 730.660 1.400 731.500 571.200 ;
    RECT 731.780 1.400 732.620 571.200 ;
    RECT 732.900 1.400 733.740 571.200 ;
    RECT 734.020 1.400 734.860 571.200 ;
    RECT 735.140 1.400 735.980 571.200 ;
    RECT 736.260 1.400 737.100 571.200 ;
    RECT 737.380 1.400 738.220 571.200 ;
    RECT 738.500 1.400 739.340 571.200 ;
    RECT 739.620 1.400 740.460 571.200 ;
    RECT 740.740 1.400 741.580 571.200 ;
    RECT 741.860 1.400 742.700 571.200 ;
    RECT 742.980 1.400 743.820 571.200 ;
    RECT 744.100 1.400 744.940 571.200 ;
    RECT 745.220 1.400 747.080 571.200 ;
    LAYER OVERLAP ;
    RECT 0 0 747.080 572.600 ;
  END
END sram_96x4096_1rw

END LIBRARY
