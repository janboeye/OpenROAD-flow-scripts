VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_15x4096_1rw
  FOREIGN sram_15x4096_1rw 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 377.910 BY 323.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END w_mask_in[14]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.125 0.070 76.195 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.085 0.070 92.155 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.725 0.070 102.795 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.045 0.070 108.115 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.365 0.070 113.435 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.685 0.070 118.755 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.005 0.070 124.075 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.645 0.070 134.715 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.285 0.070 145.355 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END rd_out[14]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.885 0.070 150.955 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.205 0.070 156.275 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.525 0.070 161.595 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.845 0.070 166.915 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.485 0.070 177.555 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.805 0.070 182.875 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.445 0.070 193.515 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.765 0.070 198.835 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.085 0.070 204.155 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.405 0.070 209.475 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.725 0.070 214.795 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.045 0.070 220.115 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.365 0.070 225.435 ;
    END
  END wd_in[14]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.645 0.070 225.715 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.965 0.070 231.035 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.285 0.070 236.355 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.605 0.070 241.675 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.925 0.070 246.995 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.245 0.070 252.315 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.565 0.070 257.635 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.885 0.070 262.955 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.205 0.070 268.275 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.525 0.070 273.595 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.845 0.070 278.915 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.165 0.070 284.235 ;
    END
  END addr_in[11]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.445 0.070 284.515 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.765 0.070 289.835 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.085 0.070 295.155 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 322.000 ;
      RECT 3.500 1.400 3.780 322.000 ;
      RECT 5.740 1.400 6.020 322.000 ;
      RECT 7.980 1.400 8.260 322.000 ;
      RECT 10.220 1.400 10.500 322.000 ;
      RECT 12.460 1.400 12.740 322.000 ;
      RECT 14.700 1.400 14.980 322.000 ;
      RECT 16.940 1.400 17.220 322.000 ;
      RECT 19.180 1.400 19.460 322.000 ;
      RECT 21.420 1.400 21.700 322.000 ;
      RECT 23.660 1.400 23.940 322.000 ;
      RECT 25.900 1.400 26.180 322.000 ;
      RECT 28.140 1.400 28.420 322.000 ;
      RECT 30.380 1.400 30.660 322.000 ;
      RECT 32.620 1.400 32.900 322.000 ;
      RECT 34.860 1.400 35.140 322.000 ;
      RECT 37.100 1.400 37.380 322.000 ;
      RECT 39.340 1.400 39.620 322.000 ;
      RECT 41.580 1.400 41.860 322.000 ;
      RECT 43.820 1.400 44.100 322.000 ;
      RECT 46.060 1.400 46.340 322.000 ;
      RECT 48.300 1.400 48.580 322.000 ;
      RECT 50.540 1.400 50.820 322.000 ;
      RECT 52.780 1.400 53.060 322.000 ;
      RECT 55.020 1.400 55.300 322.000 ;
      RECT 57.260 1.400 57.540 322.000 ;
      RECT 59.500 1.400 59.780 322.000 ;
      RECT 61.740 1.400 62.020 322.000 ;
      RECT 63.980 1.400 64.260 322.000 ;
      RECT 66.220 1.400 66.500 322.000 ;
      RECT 68.460 1.400 68.740 322.000 ;
      RECT 70.700 1.400 70.980 322.000 ;
      RECT 72.940 1.400 73.220 322.000 ;
      RECT 75.180 1.400 75.460 322.000 ;
      RECT 77.420 1.400 77.700 322.000 ;
      RECT 79.660 1.400 79.940 322.000 ;
      RECT 81.900 1.400 82.180 322.000 ;
      RECT 84.140 1.400 84.420 322.000 ;
      RECT 86.380 1.400 86.660 322.000 ;
      RECT 88.620 1.400 88.900 322.000 ;
      RECT 90.860 1.400 91.140 322.000 ;
      RECT 93.100 1.400 93.380 322.000 ;
      RECT 95.340 1.400 95.620 322.000 ;
      RECT 97.580 1.400 97.860 322.000 ;
      RECT 99.820 1.400 100.100 322.000 ;
      RECT 102.060 1.400 102.340 322.000 ;
      RECT 104.300 1.400 104.580 322.000 ;
      RECT 106.540 1.400 106.820 322.000 ;
      RECT 108.780 1.400 109.060 322.000 ;
      RECT 111.020 1.400 111.300 322.000 ;
      RECT 113.260 1.400 113.540 322.000 ;
      RECT 115.500 1.400 115.780 322.000 ;
      RECT 117.740 1.400 118.020 322.000 ;
      RECT 119.980 1.400 120.260 322.000 ;
      RECT 122.220 1.400 122.500 322.000 ;
      RECT 124.460 1.400 124.740 322.000 ;
      RECT 126.700 1.400 126.980 322.000 ;
      RECT 128.940 1.400 129.220 322.000 ;
      RECT 131.180 1.400 131.460 322.000 ;
      RECT 133.420 1.400 133.700 322.000 ;
      RECT 135.660 1.400 135.940 322.000 ;
      RECT 137.900 1.400 138.180 322.000 ;
      RECT 140.140 1.400 140.420 322.000 ;
      RECT 142.380 1.400 142.660 322.000 ;
      RECT 144.620 1.400 144.900 322.000 ;
      RECT 146.860 1.400 147.140 322.000 ;
      RECT 149.100 1.400 149.380 322.000 ;
      RECT 151.340 1.400 151.620 322.000 ;
      RECT 153.580 1.400 153.860 322.000 ;
      RECT 155.820 1.400 156.100 322.000 ;
      RECT 158.060 1.400 158.340 322.000 ;
      RECT 160.300 1.400 160.580 322.000 ;
      RECT 162.540 1.400 162.820 322.000 ;
      RECT 164.780 1.400 165.060 322.000 ;
      RECT 167.020 1.400 167.300 322.000 ;
      RECT 169.260 1.400 169.540 322.000 ;
      RECT 171.500 1.400 171.780 322.000 ;
      RECT 173.740 1.400 174.020 322.000 ;
      RECT 175.980 1.400 176.260 322.000 ;
      RECT 178.220 1.400 178.500 322.000 ;
      RECT 180.460 1.400 180.740 322.000 ;
      RECT 182.700 1.400 182.980 322.000 ;
      RECT 184.940 1.400 185.220 322.000 ;
      RECT 187.180 1.400 187.460 322.000 ;
      RECT 189.420 1.400 189.700 322.000 ;
      RECT 191.660 1.400 191.940 322.000 ;
      RECT 193.900 1.400 194.180 322.000 ;
      RECT 196.140 1.400 196.420 322.000 ;
      RECT 198.380 1.400 198.660 322.000 ;
      RECT 200.620 1.400 200.900 322.000 ;
      RECT 202.860 1.400 203.140 322.000 ;
      RECT 205.100 1.400 205.380 322.000 ;
      RECT 207.340 1.400 207.620 322.000 ;
      RECT 209.580 1.400 209.860 322.000 ;
      RECT 211.820 1.400 212.100 322.000 ;
      RECT 214.060 1.400 214.340 322.000 ;
      RECT 216.300 1.400 216.580 322.000 ;
      RECT 218.540 1.400 218.820 322.000 ;
      RECT 220.780 1.400 221.060 322.000 ;
      RECT 223.020 1.400 223.300 322.000 ;
      RECT 225.260 1.400 225.540 322.000 ;
      RECT 227.500 1.400 227.780 322.000 ;
      RECT 229.740 1.400 230.020 322.000 ;
      RECT 231.980 1.400 232.260 322.000 ;
      RECT 234.220 1.400 234.500 322.000 ;
      RECT 236.460 1.400 236.740 322.000 ;
      RECT 238.700 1.400 238.980 322.000 ;
      RECT 240.940 1.400 241.220 322.000 ;
      RECT 243.180 1.400 243.460 322.000 ;
      RECT 245.420 1.400 245.700 322.000 ;
      RECT 247.660 1.400 247.940 322.000 ;
      RECT 249.900 1.400 250.180 322.000 ;
      RECT 252.140 1.400 252.420 322.000 ;
      RECT 254.380 1.400 254.660 322.000 ;
      RECT 256.620 1.400 256.900 322.000 ;
      RECT 258.860 1.400 259.140 322.000 ;
      RECT 261.100 1.400 261.380 322.000 ;
      RECT 263.340 1.400 263.620 322.000 ;
      RECT 265.580 1.400 265.860 322.000 ;
      RECT 267.820 1.400 268.100 322.000 ;
      RECT 270.060 1.400 270.340 322.000 ;
      RECT 272.300 1.400 272.580 322.000 ;
      RECT 274.540 1.400 274.820 322.000 ;
      RECT 276.780 1.400 277.060 322.000 ;
      RECT 279.020 1.400 279.300 322.000 ;
      RECT 281.260 1.400 281.540 322.000 ;
      RECT 283.500 1.400 283.780 322.000 ;
      RECT 285.740 1.400 286.020 322.000 ;
      RECT 287.980 1.400 288.260 322.000 ;
      RECT 290.220 1.400 290.500 322.000 ;
      RECT 292.460 1.400 292.740 322.000 ;
      RECT 294.700 1.400 294.980 322.000 ;
      RECT 296.940 1.400 297.220 322.000 ;
      RECT 299.180 1.400 299.460 322.000 ;
      RECT 301.420 1.400 301.700 322.000 ;
      RECT 303.660 1.400 303.940 322.000 ;
      RECT 305.900 1.400 306.180 322.000 ;
      RECT 308.140 1.400 308.420 322.000 ;
      RECT 310.380 1.400 310.660 322.000 ;
      RECT 312.620 1.400 312.900 322.000 ;
      RECT 314.860 1.400 315.140 322.000 ;
      RECT 317.100 1.400 317.380 322.000 ;
      RECT 319.340 1.400 319.620 322.000 ;
      RECT 321.580 1.400 321.860 322.000 ;
      RECT 323.820 1.400 324.100 322.000 ;
      RECT 326.060 1.400 326.340 322.000 ;
      RECT 328.300 1.400 328.580 322.000 ;
      RECT 330.540 1.400 330.820 322.000 ;
      RECT 332.780 1.400 333.060 322.000 ;
      RECT 335.020 1.400 335.300 322.000 ;
      RECT 337.260 1.400 337.540 322.000 ;
      RECT 339.500 1.400 339.780 322.000 ;
      RECT 341.740 1.400 342.020 322.000 ;
      RECT 343.980 1.400 344.260 322.000 ;
      RECT 346.220 1.400 346.500 322.000 ;
      RECT 348.460 1.400 348.740 322.000 ;
      RECT 350.700 1.400 350.980 322.000 ;
      RECT 352.940 1.400 353.220 322.000 ;
      RECT 355.180 1.400 355.460 322.000 ;
      RECT 357.420 1.400 357.700 322.000 ;
      RECT 359.660 1.400 359.940 322.000 ;
      RECT 361.900 1.400 362.180 322.000 ;
      RECT 364.140 1.400 364.420 322.000 ;
      RECT 366.380 1.400 366.660 322.000 ;
      RECT 368.620 1.400 368.900 322.000 ;
      RECT 370.860 1.400 371.140 322.000 ;
      RECT 373.100 1.400 373.380 322.000 ;
      RECT 375.340 1.400 375.620 322.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 322.000 ;
      RECT 4.620 1.400 4.900 322.000 ;
      RECT 6.860 1.400 7.140 322.000 ;
      RECT 9.100 1.400 9.380 322.000 ;
      RECT 11.340 1.400 11.620 322.000 ;
      RECT 13.580 1.400 13.860 322.000 ;
      RECT 15.820 1.400 16.100 322.000 ;
      RECT 18.060 1.400 18.340 322.000 ;
      RECT 20.300 1.400 20.580 322.000 ;
      RECT 22.540 1.400 22.820 322.000 ;
      RECT 24.780 1.400 25.060 322.000 ;
      RECT 27.020 1.400 27.300 322.000 ;
      RECT 29.260 1.400 29.540 322.000 ;
      RECT 31.500 1.400 31.780 322.000 ;
      RECT 33.740 1.400 34.020 322.000 ;
      RECT 35.980 1.400 36.260 322.000 ;
      RECT 38.220 1.400 38.500 322.000 ;
      RECT 40.460 1.400 40.740 322.000 ;
      RECT 42.700 1.400 42.980 322.000 ;
      RECT 44.940 1.400 45.220 322.000 ;
      RECT 47.180 1.400 47.460 322.000 ;
      RECT 49.420 1.400 49.700 322.000 ;
      RECT 51.660 1.400 51.940 322.000 ;
      RECT 53.900 1.400 54.180 322.000 ;
      RECT 56.140 1.400 56.420 322.000 ;
      RECT 58.380 1.400 58.660 322.000 ;
      RECT 60.620 1.400 60.900 322.000 ;
      RECT 62.860 1.400 63.140 322.000 ;
      RECT 65.100 1.400 65.380 322.000 ;
      RECT 67.340 1.400 67.620 322.000 ;
      RECT 69.580 1.400 69.860 322.000 ;
      RECT 71.820 1.400 72.100 322.000 ;
      RECT 74.060 1.400 74.340 322.000 ;
      RECT 76.300 1.400 76.580 322.000 ;
      RECT 78.540 1.400 78.820 322.000 ;
      RECT 80.780 1.400 81.060 322.000 ;
      RECT 83.020 1.400 83.300 322.000 ;
      RECT 85.260 1.400 85.540 322.000 ;
      RECT 87.500 1.400 87.780 322.000 ;
      RECT 89.740 1.400 90.020 322.000 ;
      RECT 91.980 1.400 92.260 322.000 ;
      RECT 94.220 1.400 94.500 322.000 ;
      RECT 96.460 1.400 96.740 322.000 ;
      RECT 98.700 1.400 98.980 322.000 ;
      RECT 100.940 1.400 101.220 322.000 ;
      RECT 103.180 1.400 103.460 322.000 ;
      RECT 105.420 1.400 105.700 322.000 ;
      RECT 107.660 1.400 107.940 322.000 ;
      RECT 109.900 1.400 110.180 322.000 ;
      RECT 112.140 1.400 112.420 322.000 ;
      RECT 114.380 1.400 114.660 322.000 ;
      RECT 116.620 1.400 116.900 322.000 ;
      RECT 118.860 1.400 119.140 322.000 ;
      RECT 121.100 1.400 121.380 322.000 ;
      RECT 123.340 1.400 123.620 322.000 ;
      RECT 125.580 1.400 125.860 322.000 ;
      RECT 127.820 1.400 128.100 322.000 ;
      RECT 130.060 1.400 130.340 322.000 ;
      RECT 132.300 1.400 132.580 322.000 ;
      RECT 134.540 1.400 134.820 322.000 ;
      RECT 136.780 1.400 137.060 322.000 ;
      RECT 139.020 1.400 139.300 322.000 ;
      RECT 141.260 1.400 141.540 322.000 ;
      RECT 143.500 1.400 143.780 322.000 ;
      RECT 145.740 1.400 146.020 322.000 ;
      RECT 147.980 1.400 148.260 322.000 ;
      RECT 150.220 1.400 150.500 322.000 ;
      RECT 152.460 1.400 152.740 322.000 ;
      RECT 154.700 1.400 154.980 322.000 ;
      RECT 156.940 1.400 157.220 322.000 ;
      RECT 159.180 1.400 159.460 322.000 ;
      RECT 161.420 1.400 161.700 322.000 ;
      RECT 163.660 1.400 163.940 322.000 ;
      RECT 165.900 1.400 166.180 322.000 ;
      RECT 168.140 1.400 168.420 322.000 ;
      RECT 170.380 1.400 170.660 322.000 ;
      RECT 172.620 1.400 172.900 322.000 ;
      RECT 174.860 1.400 175.140 322.000 ;
      RECT 177.100 1.400 177.380 322.000 ;
      RECT 179.340 1.400 179.620 322.000 ;
      RECT 181.580 1.400 181.860 322.000 ;
      RECT 183.820 1.400 184.100 322.000 ;
      RECT 186.060 1.400 186.340 322.000 ;
      RECT 188.300 1.400 188.580 322.000 ;
      RECT 190.540 1.400 190.820 322.000 ;
      RECT 192.780 1.400 193.060 322.000 ;
      RECT 195.020 1.400 195.300 322.000 ;
      RECT 197.260 1.400 197.540 322.000 ;
      RECT 199.500 1.400 199.780 322.000 ;
      RECT 201.740 1.400 202.020 322.000 ;
      RECT 203.980 1.400 204.260 322.000 ;
      RECT 206.220 1.400 206.500 322.000 ;
      RECT 208.460 1.400 208.740 322.000 ;
      RECT 210.700 1.400 210.980 322.000 ;
      RECT 212.940 1.400 213.220 322.000 ;
      RECT 215.180 1.400 215.460 322.000 ;
      RECT 217.420 1.400 217.700 322.000 ;
      RECT 219.660 1.400 219.940 322.000 ;
      RECT 221.900 1.400 222.180 322.000 ;
      RECT 224.140 1.400 224.420 322.000 ;
      RECT 226.380 1.400 226.660 322.000 ;
      RECT 228.620 1.400 228.900 322.000 ;
      RECT 230.860 1.400 231.140 322.000 ;
      RECT 233.100 1.400 233.380 322.000 ;
      RECT 235.340 1.400 235.620 322.000 ;
      RECT 237.580 1.400 237.860 322.000 ;
      RECT 239.820 1.400 240.100 322.000 ;
      RECT 242.060 1.400 242.340 322.000 ;
      RECT 244.300 1.400 244.580 322.000 ;
      RECT 246.540 1.400 246.820 322.000 ;
      RECT 248.780 1.400 249.060 322.000 ;
      RECT 251.020 1.400 251.300 322.000 ;
      RECT 253.260 1.400 253.540 322.000 ;
      RECT 255.500 1.400 255.780 322.000 ;
      RECT 257.740 1.400 258.020 322.000 ;
      RECT 259.980 1.400 260.260 322.000 ;
      RECT 262.220 1.400 262.500 322.000 ;
      RECT 264.460 1.400 264.740 322.000 ;
      RECT 266.700 1.400 266.980 322.000 ;
      RECT 268.940 1.400 269.220 322.000 ;
      RECT 271.180 1.400 271.460 322.000 ;
      RECT 273.420 1.400 273.700 322.000 ;
      RECT 275.660 1.400 275.940 322.000 ;
      RECT 277.900 1.400 278.180 322.000 ;
      RECT 280.140 1.400 280.420 322.000 ;
      RECT 282.380 1.400 282.660 322.000 ;
      RECT 284.620 1.400 284.900 322.000 ;
      RECT 286.860 1.400 287.140 322.000 ;
      RECT 289.100 1.400 289.380 322.000 ;
      RECT 291.340 1.400 291.620 322.000 ;
      RECT 293.580 1.400 293.860 322.000 ;
      RECT 295.820 1.400 296.100 322.000 ;
      RECT 298.060 1.400 298.340 322.000 ;
      RECT 300.300 1.400 300.580 322.000 ;
      RECT 302.540 1.400 302.820 322.000 ;
      RECT 304.780 1.400 305.060 322.000 ;
      RECT 307.020 1.400 307.300 322.000 ;
      RECT 309.260 1.400 309.540 322.000 ;
      RECT 311.500 1.400 311.780 322.000 ;
      RECT 313.740 1.400 314.020 322.000 ;
      RECT 315.980 1.400 316.260 322.000 ;
      RECT 318.220 1.400 318.500 322.000 ;
      RECT 320.460 1.400 320.740 322.000 ;
      RECT 322.700 1.400 322.980 322.000 ;
      RECT 324.940 1.400 325.220 322.000 ;
      RECT 327.180 1.400 327.460 322.000 ;
      RECT 329.420 1.400 329.700 322.000 ;
      RECT 331.660 1.400 331.940 322.000 ;
      RECT 333.900 1.400 334.180 322.000 ;
      RECT 336.140 1.400 336.420 322.000 ;
      RECT 338.380 1.400 338.660 322.000 ;
      RECT 340.620 1.400 340.900 322.000 ;
      RECT 342.860 1.400 343.140 322.000 ;
      RECT 345.100 1.400 345.380 322.000 ;
      RECT 347.340 1.400 347.620 322.000 ;
      RECT 349.580 1.400 349.860 322.000 ;
      RECT 351.820 1.400 352.100 322.000 ;
      RECT 354.060 1.400 354.340 322.000 ;
      RECT 356.300 1.400 356.580 322.000 ;
      RECT 358.540 1.400 358.820 322.000 ;
      RECT 360.780 1.400 361.060 322.000 ;
      RECT 363.020 1.400 363.300 322.000 ;
      RECT 365.260 1.400 365.540 322.000 ;
      RECT 367.500 1.400 367.780 322.000 ;
      RECT 369.740 1.400 370.020 322.000 ;
      RECT 371.980 1.400 372.260 322.000 ;
      RECT 374.220 1.400 374.500 322.000 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 377.910 323.400 ;
    LAYER metal2 ;
    RECT 0 0 377.910 323.400 ;
    LAYER metal3 ;
    RECT 0.070 0 377.910 323.400 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 6.685 ;
    RECT 0 6.755 0.070 12.005 ;
    RECT 0 12.075 0.070 17.325 ;
    RECT 0 17.395 0.070 22.645 ;
    RECT 0 22.715 0.070 27.965 ;
    RECT 0 28.035 0.070 33.285 ;
    RECT 0 33.355 0.070 38.605 ;
    RECT 0 38.675 0.070 43.925 ;
    RECT 0 43.995 0.070 49.245 ;
    RECT 0 49.315 0.070 54.565 ;
    RECT 0 54.635 0.070 59.885 ;
    RECT 0 59.955 0.070 65.205 ;
    RECT 0 65.275 0.070 70.525 ;
    RECT 0 70.595 0.070 75.845 ;
    RECT 0 75.915 0.070 76.125 ;
    RECT 0 76.195 0.070 81.445 ;
    RECT 0 81.515 0.070 86.765 ;
    RECT 0 86.835 0.070 92.085 ;
    RECT 0 92.155 0.070 97.405 ;
    RECT 0 97.475 0.070 102.725 ;
    RECT 0 102.795 0.070 108.045 ;
    RECT 0 108.115 0.070 113.365 ;
    RECT 0 113.435 0.070 118.685 ;
    RECT 0 118.755 0.070 124.005 ;
    RECT 0 124.075 0.070 129.325 ;
    RECT 0 129.395 0.070 134.645 ;
    RECT 0 134.715 0.070 139.965 ;
    RECT 0 140.035 0.070 145.285 ;
    RECT 0 145.355 0.070 150.605 ;
    RECT 0 150.675 0.070 150.885 ;
    RECT 0 150.955 0.070 156.205 ;
    RECT 0 156.275 0.070 161.525 ;
    RECT 0 161.595 0.070 166.845 ;
    RECT 0 166.915 0.070 172.165 ;
    RECT 0 172.235 0.070 177.485 ;
    RECT 0 177.555 0.070 182.805 ;
    RECT 0 182.875 0.070 188.125 ;
    RECT 0 188.195 0.070 193.445 ;
    RECT 0 193.515 0.070 198.765 ;
    RECT 0 198.835 0.070 204.085 ;
    RECT 0 204.155 0.070 209.405 ;
    RECT 0 209.475 0.070 214.725 ;
    RECT 0 214.795 0.070 220.045 ;
    RECT 0 220.115 0.070 225.365 ;
    RECT 0 225.435 0.070 225.645 ;
    RECT 0 225.715 0.070 230.965 ;
    RECT 0 231.035 0.070 236.285 ;
    RECT 0 236.355 0.070 241.605 ;
    RECT 0 241.675 0.070 246.925 ;
    RECT 0 246.995 0.070 252.245 ;
    RECT 0 252.315 0.070 257.565 ;
    RECT 0 257.635 0.070 262.885 ;
    RECT 0 262.955 0.070 268.205 ;
    RECT 0 268.275 0.070 273.525 ;
    RECT 0 273.595 0.070 278.845 ;
    RECT 0 278.915 0.070 284.165 ;
    RECT 0 284.235 0.070 284.445 ;
    RECT 0 284.515 0.070 289.765 ;
    RECT 0 289.835 0.070 295.085 ;
    RECT 0 295.155 0.070 323.400 ;
    LAYER metal4 ;
    RECT 0 0 377.910 1.400 ;
    RECT 0 322.000 377.910 323.400 ;
    RECT 0.000 1.400 1.260 322.000 ;
    RECT 1.540 1.400 2.380 322.000 ;
    RECT 2.660 1.400 3.500 322.000 ;
    RECT 3.780 1.400 4.620 322.000 ;
    RECT 4.900 1.400 5.740 322.000 ;
    RECT 6.020 1.400 6.860 322.000 ;
    RECT 7.140 1.400 7.980 322.000 ;
    RECT 8.260 1.400 9.100 322.000 ;
    RECT 9.380 1.400 10.220 322.000 ;
    RECT 10.500 1.400 11.340 322.000 ;
    RECT 11.620 1.400 12.460 322.000 ;
    RECT 12.740 1.400 13.580 322.000 ;
    RECT 13.860 1.400 14.700 322.000 ;
    RECT 14.980 1.400 15.820 322.000 ;
    RECT 16.100 1.400 16.940 322.000 ;
    RECT 17.220 1.400 18.060 322.000 ;
    RECT 18.340 1.400 19.180 322.000 ;
    RECT 19.460 1.400 20.300 322.000 ;
    RECT 20.580 1.400 21.420 322.000 ;
    RECT 21.700 1.400 22.540 322.000 ;
    RECT 22.820 1.400 23.660 322.000 ;
    RECT 23.940 1.400 24.780 322.000 ;
    RECT 25.060 1.400 25.900 322.000 ;
    RECT 26.180 1.400 27.020 322.000 ;
    RECT 27.300 1.400 28.140 322.000 ;
    RECT 28.420 1.400 29.260 322.000 ;
    RECT 29.540 1.400 30.380 322.000 ;
    RECT 30.660 1.400 31.500 322.000 ;
    RECT 31.780 1.400 32.620 322.000 ;
    RECT 32.900 1.400 33.740 322.000 ;
    RECT 34.020 1.400 34.860 322.000 ;
    RECT 35.140 1.400 35.980 322.000 ;
    RECT 36.260 1.400 37.100 322.000 ;
    RECT 37.380 1.400 38.220 322.000 ;
    RECT 38.500 1.400 39.340 322.000 ;
    RECT 39.620 1.400 40.460 322.000 ;
    RECT 40.740 1.400 41.580 322.000 ;
    RECT 41.860 1.400 42.700 322.000 ;
    RECT 42.980 1.400 43.820 322.000 ;
    RECT 44.100 1.400 44.940 322.000 ;
    RECT 45.220 1.400 46.060 322.000 ;
    RECT 46.340 1.400 47.180 322.000 ;
    RECT 47.460 1.400 48.300 322.000 ;
    RECT 48.580 1.400 49.420 322.000 ;
    RECT 49.700 1.400 50.540 322.000 ;
    RECT 50.820 1.400 51.660 322.000 ;
    RECT 51.940 1.400 52.780 322.000 ;
    RECT 53.060 1.400 53.900 322.000 ;
    RECT 54.180 1.400 55.020 322.000 ;
    RECT 55.300 1.400 56.140 322.000 ;
    RECT 56.420 1.400 57.260 322.000 ;
    RECT 57.540 1.400 58.380 322.000 ;
    RECT 58.660 1.400 59.500 322.000 ;
    RECT 59.780 1.400 60.620 322.000 ;
    RECT 60.900 1.400 61.740 322.000 ;
    RECT 62.020 1.400 62.860 322.000 ;
    RECT 63.140 1.400 63.980 322.000 ;
    RECT 64.260 1.400 65.100 322.000 ;
    RECT 65.380 1.400 66.220 322.000 ;
    RECT 66.500 1.400 67.340 322.000 ;
    RECT 67.620 1.400 68.460 322.000 ;
    RECT 68.740 1.400 69.580 322.000 ;
    RECT 69.860 1.400 70.700 322.000 ;
    RECT 70.980 1.400 71.820 322.000 ;
    RECT 72.100 1.400 72.940 322.000 ;
    RECT 73.220 1.400 74.060 322.000 ;
    RECT 74.340 1.400 75.180 322.000 ;
    RECT 75.460 1.400 76.300 322.000 ;
    RECT 76.580 1.400 77.420 322.000 ;
    RECT 77.700 1.400 78.540 322.000 ;
    RECT 78.820 1.400 79.660 322.000 ;
    RECT 79.940 1.400 80.780 322.000 ;
    RECT 81.060 1.400 81.900 322.000 ;
    RECT 82.180 1.400 83.020 322.000 ;
    RECT 83.300 1.400 84.140 322.000 ;
    RECT 84.420 1.400 85.260 322.000 ;
    RECT 85.540 1.400 86.380 322.000 ;
    RECT 86.660 1.400 87.500 322.000 ;
    RECT 87.780 1.400 88.620 322.000 ;
    RECT 88.900 1.400 89.740 322.000 ;
    RECT 90.020 1.400 90.860 322.000 ;
    RECT 91.140 1.400 91.980 322.000 ;
    RECT 92.260 1.400 93.100 322.000 ;
    RECT 93.380 1.400 94.220 322.000 ;
    RECT 94.500 1.400 95.340 322.000 ;
    RECT 95.620 1.400 96.460 322.000 ;
    RECT 96.740 1.400 97.580 322.000 ;
    RECT 97.860 1.400 98.700 322.000 ;
    RECT 98.980 1.400 99.820 322.000 ;
    RECT 100.100 1.400 100.940 322.000 ;
    RECT 101.220 1.400 102.060 322.000 ;
    RECT 102.340 1.400 103.180 322.000 ;
    RECT 103.460 1.400 104.300 322.000 ;
    RECT 104.580 1.400 105.420 322.000 ;
    RECT 105.700 1.400 106.540 322.000 ;
    RECT 106.820 1.400 107.660 322.000 ;
    RECT 107.940 1.400 108.780 322.000 ;
    RECT 109.060 1.400 109.900 322.000 ;
    RECT 110.180 1.400 111.020 322.000 ;
    RECT 111.300 1.400 112.140 322.000 ;
    RECT 112.420 1.400 113.260 322.000 ;
    RECT 113.540 1.400 114.380 322.000 ;
    RECT 114.660 1.400 115.500 322.000 ;
    RECT 115.780 1.400 116.620 322.000 ;
    RECT 116.900 1.400 117.740 322.000 ;
    RECT 118.020 1.400 118.860 322.000 ;
    RECT 119.140 1.400 119.980 322.000 ;
    RECT 120.260 1.400 121.100 322.000 ;
    RECT 121.380 1.400 122.220 322.000 ;
    RECT 122.500 1.400 123.340 322.000 ;
    RECT 123.620 1.400 124.460 322.000 ;
    RECT 124.740 1.400 125.580 322.000 ;
    RECT 125.860 1.400 126.700 322.000 ;
    RECT 126.980 1.400 127.820 322.000 ;
    RECT 128.100 1.400 128.940 322.000 ;
    RECT 129.220 1.400 130.060 322.000 ;
    RECT 130.340 1.400 131.180 322.000 ;
    RECT 131.460 1.400 132.300 322.000 ;
    RECT 132.580 1.400 133.420 322.000 ;
    RECT 133.700 1.400 134.540 322.000 ;
    RECT 134.820 1.400 135.660 322.000 ;
    RECT 135.940 1.400 136.780 322.000 ;
    RECT 137.060 1.400 137.900 322.000 ;
    RECT 138.180 1.400 139.020 322.000 ;
    RECT 139.300 1.400 140.140 322.000 ;
    RECT 140.420 1.400 141.260 322.000 ;
    RECT 141.540 1.400 142.380 322.000 ;
    RECT 142.660 1.400 143.500 322.000 ;
    RECT 143.780 1.400 144.620 322.000 ;
    RECT 144.900 1.400 145.740 322.000 ;
    RECT 146.020 1.400 146.860 322.000 ;
    RECT 147.140 1.400 147.980 322.000 ;
    RECT 148.260 1.400 149.100 322.000 ;
    RECT 149.380 1.400 150.220 322.000 ;
    RECT 150.500 1.400 151.340 322.000 ;
    RECT 151.620 1.400 152.460 322.000 ;
    RECT 152.740 1.400 153.580 322.000 ;
    RECT 153.860 1.400 154.700 322.000 ;
    RECT 154.980 1.400 155.820 322.000 ;
    RECT 156.100 1.400 156.940 322.000 ;
    RECT 157.220 1.400 158.060 322.000 ;
    RECT 158.340 1.400 159.180 322.000 ;
    RECT 159.460 1.400 160.300 322.000 ;
    RECT 160.580 1.400 161.420 322.000 ;
    RECT 161.700 1.400 162.540 322.000 ;
    RECT 162.820 1.400 163.660 322.000 ;
    RECT 163.940 1.400 164.780 322.000 ;
    RECT 165.060 1.400 165.900 322.000 ;
    RECT 166.180 1.400 167.020 322.000 ;
    RECT 167.300 1.400 168.140 322.000 ;
    RECT 168.420 1.400 169.260 322.000 ;
    RECT 169.540 1.400 170.380 322.000 ;
    RECT 170.660 1.400 171.500 322.000 ;
    RECT 171.780 1.400 172.620 322.000 ;
    RECT 172.900 1.400 173.740 322.000 ;
    RECT 174.020 1.400 174.860 322.000 ;
    RECT 175.140 1.400 175.980 322.000 ;
    RECT 176.260 1.400 177.100 322.000 ;
    RECT 177.380 1.400 178.220 322.000 ;
    RECT 178.500 1.400 179.340 322.000 ;
    RECT 179.620 1.400 180.460 322.000 ;
    RECT 180.740 1.400 181.580 322.000 ;
    RECT 181.860 1.400 182.700 322.000 ;
    RECT 182.980 1.400 183.820 322.000 ;
    RECT 184.100 1.400 184.940 322.000 ;
    RECT 185.220 1.400 186.060 322.000 ;
    RECT 186.340 1.400 187.180 322.000 ;
    RECT 187.460 1.400 188.300 322.000 ;
    RECT 188.580 1.400 189.420 322.000 ;
    RECT 189.700 1.400 190.540 322.000 ;
    RECT 190.820 1.400 191.660 322.000 ;
    RECT 191.940 1.400 192.780 322.000 ;
    RECT 193.060 1.400 193.900 322.000 ;
    RECT 194.180 1.400 195.020 322.000 ;
    RECT 195.300 1.400 196.140 322.000 ;
    RECT 196.420 1.400 197.260 322.000 ;
    RECT 197.540 1.400 198.380 322.000 ;
    RECT 198.660 1.400 199.500 322.000 ;
    RECT 199.780 1.400 200.620 322.000 ;
    RECT 200.900 1.400 201.740 322.000 ;
    RECT 202.020 1.400 202.860 322.000 ;
    RECT 203.140 1.400 203.980 322.000 ;
    RECT 204.260 1.400 205.100 322.000 ;
    RECT 205.380 1.400 206.220 322.000 ;
    RECT 206.500 1.400 207.340 322.000 ;
    RECT 207.620 1.400 208.460 322.000 ;
    RECT 208.740 1.400 209.580 322.000 ;
    RECT 209.860 1.400 210.700 322.000 ;
    RECT 210.980 1.400 211.820 322.000 ;
    RECT 212.100 1.400 212.940 322.000 ;
    RECT 213.220 1.400 214.060 322.000 ;
    RECT 214.340 1.400 215.180 322.000 ;
    RECT 215.460 1.400 216.300 322.000 ;
    RECT 216.580 1.400 217.420 322.000 ;
    RECT 217.700 1.400 218.540 322.000 ;
    RECT 218.820 1.400 219.660 322.000 ;
    RECT 219.940 1.400 220.780 322.000 ;
    RECT 221.060 1.400 221.900 322.000 ;
    RECT 222.180 1.400 223.020 322.000 ;
    RECT 223.300 1.400 224.140 322.000 ;
    RECT 224.420 1.400 225.260 322.000 ;
    RECT 225.540 1.400 226.380 322.000 ;
    RECT 226.660 1.400 227.500 322.000 ;
    RECT 227.780 1.400 228.620 322.000 ;
    RECT 228.900 1.400 229.740 322.000 ;
    RECT 230.020 1.400 230.860 322.000 ;
    RECT 231.140 1.400 231.980 322.000 ;
    RECT 232.260 1.400 233.100 322.000 ;
    RECT 233.380 1.400 234.220 322.000 ;
    RECT 234.500 1.400 235.340 322.000 ;
    RECT 235.620 1.400 236.460 322.000 ;
    RECT 236.740 1.400 237.580 322.000 ;
    RECT 237.860 1.400 238.700 322.000 ;
    RECT 238.980 1.400 239.820 322.000 ;
    RECT 240.100 1.400 240.940 322.000 ;
    RECT 241.220 1.400 242.060 322.000 ;
    RECT 242.340 1.400 243.180 322.000 ;
    RECT 243.460 1.400 244.300 322.000 ;
    RECT 244.580 1.400 245.420 322.000 ;
    RECT 245.700 1.400 246.540 322.000 ;
    RECT 246.820 1.400 247.660 322.000 ;
    RECT 247.940 1.400 248.780 322.000 ;
    RECT 249.060 1.400 249.900 322.000 ;
    RECT 250.180 1.400 251.020 322.000 ;
    RECT 251.300 1.400 252.140 322.000 ;
    RECT 252.420 1.400 253.260 322.000 ;
    RECT 253.540 1.400 254.380 322.000 ;
    RECT 254.660 1.400 255.500 322.000 ;
    RECT 255.780 1.400 256.620 322.000 ;
    RECT 256.900 1.400 257.740 322.000 ;
    RECT 258.020 1.400 258.860 322.000 ;
    RECT 259.140 1.400 259.980 322.000 ;
    RECT 260.260 1.400 261.100 322.000 ;
    RECT 261.380 1.400 262.220 322.000 ;
    RECT 262.500 1.400 263.340 322.000 ;
    RECT 263.620 1.400 264.460 322.000 ;
    RECT 264.740 1.400 265.580 322.000 ;
    RECT 265.860 1.400 266.700 322.000 ;
    RECT 266.980 1.400 267.820 322.000 ;
    RECT 268.100 1.400 268.940 322.000 ;
    RECT 269.220 1.400 270.060 322.000 ;
    RECT 270.340 1.400 271.180 322.000 ;
    RECT 271.460 1.400 272.300 322.000 ;
    RECT 272.580 1.400 273.420 322.000 ;
    RECT 273.700 1.400 274.540 322.000 ;
    RECT 274.820 1.400 275.660 322.000 ;
    RECT 275.940 1.400 276.780 322.000 ;
    RECT 277.060 1.400 277.900 322.000 ;
    RECT 278.180 1.400 279.020 322.000 ;
    RECT 279.300 1.400 280.140 322.000 ;
    RECT 280.420 1.400 281.260 322.000 ;
    RECT 281.540 1.400 282.380 322.000 ;
    RECT 282.660 1.400 283.500 322.000 ;
    RECT 283.780 1.400 284.620 322.000 ;
    RECT 284.900 1.400 285.740 322.000 ;
    RECT 286.020 1.400 286.860 322.000 ;
    RECT 287.140 1.400 287.980 322.000 ;
    RECT 288.260 1.400 289.100 322.000 ;
    RECT 289.380 1.400 290.220 322.000 ;
    RECT 290.500 1.400 291.340 322.000 ;
    RECT 291.620 1.400 292.460 322.000 ;
    RECT 292.740 1.400 293.580 322.000 ;
    RECT 293.860 1.400 294.700 322.000 ;
    RECT 294.980 1.400 295.820 322.000 ;
    RECT 296.100 1.400 296.940 322.000 ;
    RECT 297.220 1.400 298.060 322.000 ;
    RECT 298.340 1.400 299.180 322.000 ;
    RECT 299.460 1.400 300.300 322.000 ;
    RECT 300.580 1.400 301.420 322.000 ;
    RECT 301.700 1.400 302.540 322.000 ;
    RECT 302.820 1.400 303.660 322.000 ;
    RECT 303.940 1.400 304.780 322.000 ;
    RECT 305.060 1.400 305.900 322.000 ;
    RECT 306.180 1.400 307.020 322.000 ;
    RECT 307.300 1.400 308.140 322.000 ;
    RECT 308.420 1.400 309.260 322.000 ;
    RECT 309.540 1.400 310.380 322.000 ;
    RECT 310.660 1.400 311.500 322.000 ;
    RECT 311.780 1.400 312.620 322.000 ;
    RECT 312.900 1.400 313.740 322.000 ;
    RECT 314.020 1.400 314.860 322.000 ;
    RECT 315.140 1.400 315.980 322.000 ;
    RECT 316.260 1.400 317.100 322.000 ;
    RECT 317.380 1.400 318.220 322.000 ;
    RECT 318.500 1.400 319.340 322.000 ;
    RECT 319.620 1.400 320.460 322.000 ;
    RECT 320.740 1.400 321.580 322.000 ;
    RECT 321.860 1.400 322.700 322.000 ;
    RECT 322.980 1.400 323.820 322.000 ;
    RECT 324.100 1.400 324.940 322.000 ;
    RECT 325.220 1.400 326.060 322.000 ;
    RECT 326.340 1.400 327.180 322.000 ;
    RECT 327.460 1.400 328.300 322.000 ;
    RECT 328.580 1.400 329.420 322.000 ;
    RECT 329.700 1.400 330.540 322.000 ;
    RECT 330.820 1.400 331.660 322.000 ;
    RECT 331.940 1.400 332.780 322.000 ;
    RECT 333.060 1.400 333.900 322.000 ;
    RECT 334.180 1.400 335.020 322.000 ;
    RECT 335.300 1.400 336.140 322.000 ;
    RECT 336.420 1.400 337.260 322.000 ;
    RECT 337.540 1.400 338.380 322.000 ;
    RECT 338.660 1.400 339.500 322.000 ;
    RECT 339.780 1.400 340.620 322.000 ;
    RECT 340.900 1.400 341.740 322.000 ;
    RECT 342.020 1.400 342.860 322.000 ;
    RECT 343.140 1.400 343.980 322.000 ;
    RECT 344.260 1.400 345.100 322.000 ;
    RECT 345.380 1.400 346.220 322.000 ;
    RECT 346.500 1.400 347.340 322.000 ;
    RECT 347.620 1.400 348.460 322.000 ;
    RECT 348.740 1.400 349.580 322.000 ;
    RECT 349.860 1.400 350.700 322.000 ;
    RECT 350.980 1.400 351.820 322.000 ;
    RECT 352.100 1.400 352.940 322.000 ;
    RECT 353.220 1.400 354.060 322.000 ;
    RECT 354.340 1.400 355.180 322.000 ;
    RECT 355.460 1.400 356.300 322.000 ;
    RECT 356.580 1.400 357.420 322.000 ;
    RECT 357.700 1.400 358.540 322.000 ;
    RECT 358.820 1.400 359.660 322.000 ;
    RECT 359.940 1.400 360.780 322.000 ;
    RECT 361.060 1.400 361.900 322.000 ;
    RECT 362.180 1.400 363.020 322.000 ;
    RECT 363.300 1.400 364.140 322.000 ;
    RECT 364.420 1.400 365.260 322.000 ;
    RECT 365.540 1.400 366.380 322.000 ;
    RECT 366.660 1.400 367.500 322.000 ;
    RECT 367.780 1.400 368.620 322.000 ;
    RECT 368.900 1.400 369.740 322.000 ;
    RECT 370.020 1.400 370.860 322.000 ;
    RECT 371.140 1.400 371.980 322.000 ;
    RECT 372.260 1.400 373.100 322.000 ;
    RECT 373.380 1.400 374.220 322.000 ;
    RECT 374.500 1.400 375.340 322.000 ;
    RECT 375.620 1.400 377.910 322.000 ;
    LAYER OVERLAP ;
    RECT 0 0 377.910 323.400 ;
  END
END sram_15x4096_1rw

END LIBRARY
