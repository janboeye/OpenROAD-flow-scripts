VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_256x4096_1rw
  FOREIGN sram_256x4096_1rw 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1631.530 BY 737.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.645 0.070 15.715 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.685 0.070 20.755 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.725 0.070 25.795 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.405 0.070 27.475 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.085 0.070 50.155 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.925 0.070 50.995 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.605 0.070 52.675 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.445 0.070 53.515 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.325 0.070 59.395 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.005 0.070 61.075 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.845 0.070 61.915 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.685 0.070 62.755 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.725 0.070 67.795 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.405 0.070 69.475 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.445 0.070 74.515 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.125 0.070 76.195 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.645 0.070 78.715 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.485 0.070 79.555 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.325 0.070 80.395 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.005 0.070 82.075 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.845 0.070 82.915 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.205 0.070 86.275 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.045 0.070 87.115 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.885 0.070 87.955 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.725 0.070 88.795 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.405 0.070 90.475 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.245 0.070 91.315 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.085 0.070 92.155 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.925 0.070 92.995 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.765 0.070 93.835 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.605 0.070 94.675 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.285 0.070 96.355 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.125 0.070 97.195 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.965 0.070 98.035 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.805 0.070 98.875 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.485 0.070 100.555 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.165 0.070 102.235 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.005 0.070 103.075 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.845 0.070 103.915 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.685 0.070 104.755 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.525 0.070 105.595 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.365 0.070 106.435 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.045 0.070 108.115 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.885 0.070 108.955 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.725 0.070 109.795 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.565 0.070 110.635 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.405 0.070 111.475 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.925 0.070 113.995 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.765 0.070 114.835 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.605 0.070 115.675 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.445 0.070 116.515 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.285 0.070 117.355 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.645 0.070 120.715 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END w_mask_in[143]
  PIN w_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.325 0.070 122.395 ;
    END
  END w_mask_in[144]
  PIN w_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.165 0.070 123.235 ;
    END
  END w_mask_in[145]
  PIN w_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.005 0.070 124.075 ;
    END
  END w_mask_in[146]
  PIN w_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END w_mask_in[147]
  PIN w_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.685 0.070 125.755 ;
    END
  END w_mask_in[148]
  PIN w_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.525 0.070 126.595 ;
    END
  END w_mask_in[149]
  PIN w_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.365 0.070 127.435 ;
    END
  END w_mask_in[150]
  PIN w_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.205 0.070 128.275 ;
    END
  END w_mask_in[151]
  PIN w_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.045 0.070 129.115 ;
    END
  END w_mask_in[152]
  PIN w_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END w_mask_in[153]
  PIN w_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END w_mask_in[154]
  PIN w_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.565 0.070 131.635 ;
    END
  END w_mask_in[155]
  PIN w_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.405 0.070 132.475 ;
    END
  END w_mask_in[156]
  PIN w_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.245 0.070 133.315 ;
    END
  END w_mask_in[157]
  PIN w_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.085 0.070 134.155 ;
    END
  END w_mask_in[158]
  PIN w_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END w_mask_in[159]
  PIN w_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.765 0.070 135.835 ;
    END
  END w_mask_in[160]
  PIN w_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END w_mask_in[161]
  PIN w_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.445 0.070 137.515 ;
    END
  END w_mask_in[162]
  PIN w_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END w_mask_in[163]
  PIN w_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END w_mask_in[164]
  PIN w_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END w_mask_in[165]
  PIN w_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.805 0.070 140.875 ;
    END
  END w_mask_in[166]
  PIN w_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END w_mask_in[167]
  PIN w_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END w_mask_in[168]
  PIN w_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END w_mask_in[169]
  PIN w_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.165 0.070 144.235 ;
    END
  END w_mask_in[170]
  PIN w_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END w_mask_in[171]
  PIN w_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.845 0.070 145.915 ;
    END
  END w_mask_in[172]
  PIN w_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END w_mask_in[173]
  PIN w_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.525 0.070 147.595 ;
    END
  END w_mask_in[174]
  PIN w_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END w_mask_in[175]
  PIN w_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.205 0.070 149.275 ;
    END
  END w_mask_in[176]
  PIN w_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.045 0.070 150.115 ;
    END
  END w_mask_in[177]
  PIN w_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.885 0.070 150.955 ;
    END
  END w_mask_in[178]
  PIN w_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.725 0.070 151.795 ;
    END
  END w_mask_in[179]
  PIN w_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.565 0.070 152.635 ;
    END
  END w_mask_in[180]
  PIN w_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.405 0.070 153.475 ;
    END
  END w_mask_in[181]
  PIN w_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END w_mask_in[182]
  PIN w_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.085 0.070 155.155 ;
    END
  END w_mask_in[183]
  PIN w_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.925 0.070 155.995 ;
    END
  END w_mask_in[184]
  PIN w_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.765 0.070 156.835 ;
    END
  END w_mask_in[185]
  PIN w_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.605 0.070 157.675 ;
    END
  END w_mask_in[186]
  PIN w_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.445 0.070 158.515 ;
    END
  END w_mask_in[187]
  PIN w_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.285 0.070 159.355 ;
    END
  END w_mask_in[188]
  PIN w_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END w_mask_in[189]
  PIN w_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.965 0.070 161.035 ;
    END
  END w_mask_in[190]
  PIN w_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.805 0.070 161.875 ;
    END
  END w_mask_in[191]
  PIN w_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.645 0.070 162.715 ;
    END
  END w_mask_in[192]
  PIN w_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.485 0.070 163.555 ;
    END
  END w_mask_in[193]
  PIN w_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.325 0.070 164.395 ;
    END
  END w_mask_in[194]
  PIN w_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END w_mask_in[195]
  PIN w_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.005 0.070 166.075 ;
    END
  END w_mask_in[196]
  PIN w_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.845 0.070 166.915 ;
    END
  END w_mask_in[197]
  PIN w_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END w_mask_in[198]
  PIN w_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.525 0.070 168.595 ;
    END
  END w_mask_in[199]
  PIN w_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.365 0.070 169.435 ;
    END
  END w_mask_in[200]
  PIN w_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END w_mask_in[201]
  PIN w_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.045 0.070 171.115 ;
    END
  END w_mask_in[202]
  PIN w_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END w_mask_in[203]
  PIN w_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.725 0.070 172.795 ;
    END
  END w_mask_in[204]
  PIN w_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.565 0.070 173.635 ;
    END
  END w_mask_in[205]
  PIN w_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.405 0.070 174.475 ;
    END
  END w_mask_in[206]
  PIN w_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.245 0.070 175.315 ;
    END
  END w_mask_in[207]
  PIN w_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.085 0.070 176.155 ;
    END
  END w_mask_in[208]
  PIN w_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.925 0.070 176.995 ;
    END
  END w_mask_in[209]
  PIN w_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END w_mask_in[210]
  PIN w_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.605 0.070 178.675 ;
    END
  END w_mask_in[211]
  PIN w_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.445 0.070 179.515 ;
    END
  END w_mask_in[212]
  PIN w_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.285 0.070 180.355 ;
    END
  END w_mask_in[213]
  PIN w_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.125 0.070 181.195 ;
    END
  END w_mask_in[214]
  PIN w_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.965 0.070 182.035 ;
    END
  END w_mask_in[215]
  PIN w_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.805 0.070 182.875 ;
    END
  END w_mask_in[216]
  PIN w_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.645 0.070 183.715 ;
    END
  END w_mask_in[217]
  PIN w_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.485 0.070 184.555 ;
    END
  END w_mask_in[218]
  PIN w_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.325 0.070 185.395 ;
    END
  END w_mask_in[219]
  PIN w_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.165 0.070 186.235 ;
    END
  END w_mask_in[220]
  PIN w_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.005 0.070 187.075 ;
    END
  END w_mask_in[221]
  PIN w_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.845 0.070 187.915 ;
    END
  END w_mask_in[222]
  PIN w_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.685 0.070 188.755 ;
    END
  END w_mask_in[223]
  PIN w_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.525 0.070 189.595 ;
    END
  END w_mask_in[224]
  PIN w_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.365 0.070 190.435 ;
    END
  END w_mask_in[225]
  PIN w_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.205 0.070 191.275 ;
    END
  END w_mask_in[226]
  PIN w_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.045 0.070 192.115 ;
    END
  END w_mask_in[227]
  PIN w_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.885 0.070 192.955 ;
    END
  END w_mask_in[228]
  PIN w_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.725 0.070 193.795 ;
    END
  END w_mask_in[229]
  PIN w_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.565 0.070 194.635 ;
    END
  END w_mask_in[230]
  PIN w_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.405 0.070 195.475 ;
    END
  END w_mask_in[231]
  PIN w_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.245 0.070 196.315 ;
    END
  END w_mask_in[232]
  PIN w_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.085 0.070 197.155 ;
    END
  END w_mask_in[233]
  PIN w_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.925 0.070 197.995 ;
    END
  END w_mask_in[234]
  PIN w_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.765 0.070 198.835 ;
    END
  END w_mask_in[235]
  PIN w_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.605 0.070 199.675 ;
    END
  END w_mask_in[236]
  PIN w_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.445 0.070 200.515 ;
    END
  END w_mask_in[237]
  PIN w_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.285 0.070 201.355 ;
    END
  END w_mask_in[238]
  PIN w_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.125 0.070 202.195 ;
    END
  END w_mask_in[239]
  PIN w_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.965 0.070 203.035 ;
    END
  END w_mask_in[240]
  PIN w_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.805 0.070 203.875 ;
    END
  END w_mask_in[241]
  PIN w_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.645 0.070 204.715 ;
    END
  END w_mask_in[242]
  PIN w_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.485 0.070 205.555 ;
    END
  END w_mask_in[243]
  PIN w_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.325 0.070 206.395 ;
    END
  END w_mask_in[244]
  PIN w_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.165 0.070 207.235 ;
    END
  END w_mask_in[245]
  PIN w_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.005 0.070 208.075 ;
    END
  END w_mask_in[246]
  PIN w_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.845 0.070 208.915 ;
    END
  END w_mask_in[247]
  PIN w_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.685 0.070 209.755 ;
    END
  END w_mask_in[248]
  PIN w_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END w_mask_in[249]
  PIN w_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.365 0.070 211.435 ;
    END
  END w_mask_in[250]
  PIN w_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.205 0.070 212.275 ;
    END
  END w_mask_in[251]
  PIN w_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.045 0.070 213.115 ;
    END
  END w_mask_in[252]
  PIN w_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.885 0.070 213.955 ;
    END
  END w_mask_in[253]
  PIN w_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.725 0.070 214.795 ;
    END
  END w_mask_in[254]
  PIN w_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.565 0.070 215.635 ;
    END
  END w_mask_in[255]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.745 0.070 234.815 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.585 0.070 235.655 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.425 0.070 236.495 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.265 0.070 237.335 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.105 0.070 238.175 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.945 0.070 239.015 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.785 0.070 239.855 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.625 0.070 240.695 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.465 0.070 241.535 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.305 0.070 242.375 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.145 0.070 243.215 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.985 0.070 244.055 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.825 0.070 244.895 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.665 0.070 245.735 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.505 0.070 246.575 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.345 0.070 247.415 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.185 0.070 248.255 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.025 0.070 249.095 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.865 0.070 249.935 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.705 0.070 250.775 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.545 0.070 251.615 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.385 0.070 252.455 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.225 0.070 253.295 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.065 0.070 254.135 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.905 0.070 254.975 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.745 0.070 255.815 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.585 0.070 256.655 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.425 0.070 257.495 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.265 0.070 258.335 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.105 0.070 259.175 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.945 0.070 260.015 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.785 0.070 260.855 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.625 0.070 261.695 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.465 0.070 262.535 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.305 0.070 263.375 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.145 0.070 264.215 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.985 0.070 265.055 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.825 0.070 265.895 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.665 0.070 266.735 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.505 0.070 267.575 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.345 0.070 268.415 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.185 0.070 269.255 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.025 0.070 270.095 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.865 0.070 270.935 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.705 0.070 271.775 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.545 0.070 272.615 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.385 0.070 273.455 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.225 0.070 274.295 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.065 0.070 275.135 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.905 0.070 275.975 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.745 0.070 276.815 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.585 0.070 277.655 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.425 0.070 278.495 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.265 0.070 279.335 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.105 0.070 280.175 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.945 0.070 281.015 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.785 0.070 281.855 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.625 0.070 282.695 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.465 0.070 283.535 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.305 0.070 284.375 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.145 0.070 285.215 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.985 0.070 286.055 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.825 0.070 286.895 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.665 0.070 287.735 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.505 0.070 288.575 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.345 0.070 289.415 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.185 0.070 290.255 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.025 0.070 291.095 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.865 0.070 291.935 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.705 0.070 292.775 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.545 0.070 293.615 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.385 0.070 294.455 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.225 0.070 295.295 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.065 0.070 296.135 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.905 0.070 296.975 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.745 0.070 297.815 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.585 0.070 298.655 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.425 0.070 299.495 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.265 0.070 300.335 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.105 0.070 301.175 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.945 0.070 302.015 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.785 0.070 302.855 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.625 0.070 303.695 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.465 0.070 304.535 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.305 0.070 305.375 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.145 0.070 306.215 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.985 0.070 307.055 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.825 0.070 307.895 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.665 0.070 308.735 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.505 0.070 309.575 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.345 0.070 310.415 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.185 0.070 311.255 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.025 0.070 312.095 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.865 0.070 312.935 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.705 0.070 313.775 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.545 0.070 314.615 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.385 0.070 315.455 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.225 0.070 316.295 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.065 0.070 317.135 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.905 0.070 317.975 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.745 0.070 318.815 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.585 0.070 319.655 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.425 0.070 320.495 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.265 0.070 321.335 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.105 0.070 322.175 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.945 0.070 323.015 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.785 0.070 323.855 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.625 0.070 324.695 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.465 0.070 325.535 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.305 0.070 326.375 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.145 0.070 327.215 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.985 0.070 328.055 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.825 0.070 328.895 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.665 0.070 329.735 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.505 0.070 330.575 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.345 0.070 331.415 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.185 0.070 332.255 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.025 0.070 333.095 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.865 0.070 333.935 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.705 0.070 334.775 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.545 0.070 335.615 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.385 0.070 336.455 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.225 0.070 337.295 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.065 0.070 338.135 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.905 0.070 338.975 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.745 0.070 339.815 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.585 0.070 340.655 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.425 0.070 341.495 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.265 0.070 342.335 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.105 0.070 343.175 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.945 0.070 344.015 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.785 0.070 344.855 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.625 0.070 345.695 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.465 0.070 346.535 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.305 0.070 347.375 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.145 0.070 348.215 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.985 0.070 349.055 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.825 0.070 349.895 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.665 0.070 350.735 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.505 0.070 351.575 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.345 0.070 352.415 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.185 0.070 353.255 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.025 0.070 354.095 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.865 0.070 354.935 ;
    END
  END rd_out[143]
  PIN rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.705 0.070 355.775 ;
    END
  END rd_out[144]
  PIN rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.545 0.070 356.615 ;
    END
  END rd_out[145]
  PIN rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.385 0.070 357.455 ;
    END
  END rd_out[146]
  PIN rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.225 0.070 358.295 ;
    END
  END rd_out[147]
  PIN rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.065 0.070 359.135 ;
    END
  END rd_out[148]
  PIN rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.905 0.070 359.975 ;
    END
  END rd_out[149]
  PIN rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.745 0.070 360.815 ;
    END
  END rd_out[150]
  PIN rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.585 0.070 361.655 ;
    END
  END rd_out[151]
  PIN rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.425 0.070 362.495 ;
    END
  END rd_out[152]
  PIN rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.265 0.070 363.335 ;
    END
  END rd_out[153]
  PIN rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.105 0.070 364.175 ;
    END
  END rd_out[154]
  PIN rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.945 0.070 365.015 ;
    END
  END rd_out[155]
  PIN rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.785 0.070 365.855 ;
    END
  END rd_out[156]
  PIN rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.625 0.070 366.695 ;
    END
  END rd_out[157]
  PIN rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.465 0.070 367.535 ;
    END
  END rd_out[158]
  PIN rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.305 0.070 368.375 ;
    END
  END rd_out[159]
  PIN rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.145 0.070 369.215 ;
    END
  END rd_out[160]
  PIN rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.985 0.070 370.055 ;
    END
  END rd_out[161]
  PIN rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.825 0.070 370.895 ;
    END
  END rd_out[162]
  PIN rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.665 0.070 371.735 ;
    END
  END rd_out[163]
  PIN rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.505 0.070 372.575 ;
    END
  END rd_out[164]
  PIN rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.345 0.070 373.415 ;
    END
  END rd_out[165]
  PIN rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.185 0.070 374.255 ;
    END
  END rd_out[166]
  PIN rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.025 0.070 375.095 ;
    END
  END rd_out[167]
  PIN rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.865 0.070 375.935 ;
    END
  END rd_out[168]
  PIN rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.705 0.070 376.775 ;
    END
  END rd_out[169]
  PIN rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.545 0.070 377.615 ;
    END
  END rd_out[170]
  PIN rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.385 0.070 378.455 ;
    END
  END rd_out[171]
  PIN rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.225 0.070 379.295 ;
    END
  END rd_out[172]
  PIN rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.065 0.070 380.135 ;
    END
  END rd_out[173]
  PIN rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.905 0.070 380.975 ;
    END
  END rd_out[174]
  PIN rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.745 0.070 381.815 ;
    END
  END rd_out[175]
  PIN rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.585 0.070 382.655 ;
    END
  END rd_out[176]
  PIN rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.425 0.070 383.495 ;
    END
  END rd_out[177]
  PIN rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.265 0.070 384.335 ;
    END
  END rd_out[178]
  PIN rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.105 0.070 385.175 ;
    END
  END rd_out[179]
  PIN rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.945 0.070 386.015 ;
    END
  END rd_out[180]
  PIN rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.785 0.070 386.855 ;
    END
  END rd_out[181]
  PIN rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.625 0.070 387.695 ;
    END
  END rd_out[182]
  PIN rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.465 0.070 388.535 ;
    END
  END rd_out[183]
  PIN rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.305 0.070 389.375 ;
    END
  END rd_out[184]
  PIN rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.145 0.070 390.215 ;
    END
  END rd_out[185]
  PIN rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.985 0.070 391.055 ;
    END
  END rd_out[186]
  PIN rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.825 0.070 391.895 ;
    END
  END rd_out[187]
  PIN rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.665 0.070 392.735 ;
    END
  END rd_out[188]
  PIN rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.505 0.070 393.575 ;
    END
  END rd_out[189]
  PIN rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.345 0.070 394.415 ;
    END
  END rd_out[190]
  PIN rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.185 0.070 395.255 ;
    END
  END rd_out[191]
  PIN rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.025 0.070 396.095 ;
    END
  END rd_out[192]
  PIN rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.865 0.070 396.935 ;
    END
  END rd_out[193]
  PIN rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.705 0.070 397.775 ;
    END
  END rd_out[194]
  PIN rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.545 0.070 398.615 ;
    END
  END rd_out[195]
  PIN rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.385 0.070 399.455 ;
    END
  END rd_out[196]
  PIN rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 400.225 0.070 400.295 ;
    END
  END rd_out[197]
  PIN rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 401.065 0.070 401.135 ;
    END
  END rd_out[198]
  PIN rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 401.905 0.070 401.975 ;
    END
  END rd_out[199]
  PIN rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 402.745 0.070 402.815 ;
    END
  END rd_out[200]
  PIN rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 403.585 0.070 403.655 ;
    END
  END rd_out[201]
  PIN rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 404.425 0.070 404.495 ;
    END
  END rd_out[202]
  PIN rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 405.265 0.070 405.335 ;
    END
  END rd_out[203]
  PIN rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 406.105 0.070 406.175 ;
    END
  END rd_out[204]
  PIN rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 406.945 0.070 407.015 ;
    END
  END rd_out[205]
  PIN rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.785 0.070 407.855 ;
    END
  END rd_out[206]
  PIN rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 408.625 0.070 408.695 ;
    END
  END rd_out[207]
  PIN rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 409.465 0.070 409.535 ;
    END
  END rd_out[208]
  PIN rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.305 0.070 410.375 ;
    END
  END rd_out[209]
  PIN rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.145 0.070 411.215 ;
    END
  END rd_out[210]
  PIN rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.985 0.070 412.055 ;
    END
  END rd_out[211]
  PIN rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 412.825 0.070 412.895 ;
    END
  END rd_out[212]
  PIN rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 413.665 0.070 413.735 ;
    END
  END rd_out[213]
  PIN rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.505 0.070 414.575 ;
    END
  END rd_out[214]
  PIN rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 415.345 0.070 415.415 ;
    END
  END rd_out[215]
  PIN rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.185 0.070 416.255 ;
    END
  END rd_out[216]
  PIN rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 417.025 0.070 417.095 ;
    END
  END rd_out[217]
  PIN rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 417.865 0.070 417.935 ;
    END
  END rd_out[218]
  PIN rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.705 0.070 418.775 ;
    END
  END rd_out[219]
  PIN rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.545 0.070 419.615 ;
    END
  END rd_out[220]
  PIN rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 420.385 0.070 420.455 ;
    END
  END rd_out[221]
  PIN rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.225 0.070 421.295 ;
    END
  END rd_out[222]
  PIN rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 422.065 0.070 422.135 ;
    END
  END rd_out[223]
  PIN rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 422.905 0.070 422.975 ;
    END
  END rd_out[224]
  PIN rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.745 0.070 423.815 ;
    END
  END rd_out[225]
  PIN rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 424.585 0.070 424.655 ;
    END
  END rd_out[226]
  PIN rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.425 0.070 425.495 ;
    END
  END rd_out[227]
  PIN rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 426.265 0.070 426.335 ;
    END
  END rd_out[228]
  PIN rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.105 0.070 427.175 ;
    END
  END rd_out[229]
  PIN rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.945 0.070 428.015 ;
    END
  END rd_out[230]
  PIN rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.785 0.070 428.855 ;
    END
  END rd_out[231]
  PIN rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 429.625 0.070 429.695 ;
    END
  END rd_out[232]
  PIN rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.465 0.070 430.535 ;
    END
  END rd_out[233]
  PIN rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 431.305 0.070 431.375 ;
    END
  END rd_out[234]
  PIN rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.145 0.070 432.215 ;
    END
  END rd_out[235]
  PIN rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.985 0.070 433.055 ;
    END
  END rd_out[236]
  PIN rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 433.825 0.070 433.895 ;
    END
  END rd_out[237]
  PIN rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 434.665 0.070 434.735 ;
    END
  END rd_out[238]
  PIN rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 435.505 0.070 435.575 ;
    END
  END rd_out[239]
  PIN rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.345 0.070 436.415 ;
    END
  END rd_out[240]
  PIN rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.185 0.070 437.255 ;
    END
  END rd_out[241]
  PIN rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.025 0.070 438.095 ;
    END
  END rd_out[242]
  PIN rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.865 0.070 438.935 ;
    END
  END rd_out[243]
  PIN rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.705 0.070 439.775 ;
    END
  END rd_out[244]
  PIN rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 440.545 0.070 440.615 ;
    END
  END rd_out[245]
  PIN rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 441.385 0.070 441.455 ;
    END
  END rd_out[246]
  PIN rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.225 0.070 442.295 ;
    END
  END rd_out[247]
  PIN rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.065 0.070 443.135 ;
    END
  END rd_out[248]
  PIN rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.905 0.070 443.975 ;
    END
  END rd_out[249]
  PIN rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.745 0.070 444.815 ;
    END
  END rd_out[250]
  PIN rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 445.585 0.070 445.655 ;
    END
  END rd_out[251]
  PIN rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.425 0.070 446.495 ;
    END
  END rd_out[252]
  PIN rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 447.265 0.070 447.335 ;
    END
  END rd_out[253]
  PIN rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.105 0.070 448.175 ;
    END
  END rd_out[254]
  PIN rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.945 0.070 449.015 ;
    END
  END rd_out[255]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.125 0.070 468.195 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.965 0.070 469.035 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 469.805 0.070 469.875 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.645 0.070 470.715 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 471.485 0.070 471.555 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.325 0.070 472.395 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 473.165 0.070 473.235 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.005 0.070 474.075 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.845 0.070 474.915 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.685 0.070 475.755 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.525 0.070 476.595 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 477.365 0.070 477.435 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 478.205 0.070 478.275 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.045 0.070 479.115 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.885 0.070 479.955 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 480.725 0.070 480.795 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.565 0.070 481.635 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 482.405 0.070 482.475 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 483.245 0.070 483.315 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.085 0.070 484.155 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.925 0.070 484.995 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 485.765 0.070 485.835 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.605 0.070 486.675 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 487.445 0.070 487.515 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 488.285 0.070 488.355 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 489.125 0.070 489.195 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 489.965 0.070 490.035 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 490.805 0.070 490.875 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 491.645 0.070 491.715 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 492.485 0.070 492.555 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.325 0.070 493.395 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 494.165 0.070 494.235 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 495.005 0.070 495.075 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 495.845 0.070 495.915 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 496.685 0.070 496.755 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 497.525 0.070 497.595 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 498.365 0.070 498.435 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 499.205 0.070 499.275 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 500.045 0.070 500.115 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 500.885 0.070 500.955 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 501.725 0.070 501.795 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 502.565 0.070 502.635 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 503.405 0.070 503.475 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.245 0.070 504.315 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.085 0.070 505.155 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.925 0.070 505.995 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.765 0.070 506.835 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.605 0.070 507.675 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.445 0.070 508.515 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.285 0.070 509.355 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.125 0.070 510.195 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.965 0.070 511.035 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.805 0.070 511.875 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.645 0.070 512.715 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.485 0.070 513.555 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.325 0.070 514.395 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.165 0.070 515.235 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.005 0.070 516.075 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.845 0.070 516.915 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.685 0.070 517.755 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.525 0.070 518.595 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.365 0.070 519.435 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.205 0.070 520.275 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.045 0.070 521.115 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.885 0.070 521.955 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.725 0.070 522.795 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.565 0.070 523.635 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.405 0.070 524.475 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.245 0.070 525.315 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.085 0.070 526.155 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.925 0.070 526.995 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.765 0.070 527.835 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.605 0.070 528.675 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.445 0.070 529.515 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.285 0.070 530.355 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.125 0.070 531.195 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.965 0.070 532.035 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.805 0.070 532.875 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.645 0.070 533.715 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.485 0.070 534.555 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.325 0.070 535.395 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.165 0.070 536.235 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.005 0.070 537.075 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.845 0.070 537.915 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.685 0.070 538.755 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.525 0.070 539.595 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.365 0.070 540.435 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.205 0.070 541.275 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.045 0.070 542.115 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.885 0.070 542.955 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.725 0.070 543.795 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.565 0.070 544.635 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.405 0.070 545.475 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.245 0.070 546.315 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.085 0.070 547.155 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.925 0.070 547.995 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.765 0.070 548.835 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.605 0.070 549.675 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.445 0.070 550.515 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.285 0.070 551.355 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.125 0.070 552.195 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.965 0.070 553.035 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.805 0.070 553.875 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.645 0.070 554.715 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.485 0.070 555.555 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.325 0.070 556.395 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.165 0.070 557.235 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.005 0.070 558.075 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.845 0.070 558.915 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.685 0.070 559.755 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.525 0.070 560.595 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.365 0.070 561.435 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.205 0.070 562.275 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.045 0.070 563.115 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.885 0.070 563.955 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.725 0.070 564.795 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.565 0.070 565.635 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.405 0.070 566.475 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.245 0.070 567.315 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.085 0.070 568.155 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.925 0.070 568.995 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.765 0.070 569.835 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.605 0.070 570.675 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.445 0.070 571.515 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.285 0.070 572.355 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.125 0.070 573.195 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.965 0.070 574.035 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.805 0.070 574.875 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.645 0.070 575.715 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.485 0.070 576.555 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.325 0.070 577.395 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.165 0.070 578.235 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.005 0.070 579.075 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.845 0.070 579.915 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.685 0.070 580.755 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.525 0.070 581.595 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.365 0.070 582.435 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.205 0.070 583.275 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.045 0.070 584.115 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.885 0.070 584.955 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.725 0.070 585.795 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.565 0.070 586.635 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.405 0.070 587.475 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.245 0.070 588.315 ;
    END
  END wd_in[143]
  PIN wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.085 0.070 589.155 ;
    END
  END wd_in[144]
  PIN wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.925 0.070 589.995 ;
    END
  END wd_in[145]
  PIN wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.765 0.070 590.835 ;
    END
  END wd_in[146]
  PIN wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.605 0.070 591.675 ;
    END
  END wd_in[147]
  PIN wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.445 0.070 592.515 ;
    END
  END wd_in[148]
  PIN wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.285 0.070 593.355 ;
    END
  END wd_in[149]
  PIN wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.125 0.070 594.195 ;
    END
  END wd_in[150]
  PIN wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.965 0.070 595.035 ;
    END
  END wd_in[151]
  PIN wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.805 0.070 595.875 ;
    END
  END wd_in[152]
  PIN wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.645 0.070 596.715 ;
    END
  END wd_in[153]
  PIN wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.485 0.070 597.555 ;
    END
  END wd_in[154]
  PIN wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.325 0.070 598.395 ;
    END
  END wd_in[155]
  PIN wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.165 0.070 599.235 ;
    END
  END wd_in[156]
  PIN wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.005 0.070 600.075 ;
    END
  END wd_in[157]
  PIN wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.845 0.070 600.915 ;
    END
  END wd_in[158]
  PIN wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.685 0.070 601.755 ;
    END
  END wd_in[159]
  PIN wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.525 0.070 602.595 ;
    END
  END wd_in[160]
  PIN wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.365 0.070 603.435 ;
    END
  END wd_in[161]
  PIN wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.205 0.070 604.275 ;
    END
  END wd_in[162]
  PIN wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.045 0.070 605.115 ;
    END
  END wd_in[163]
  PIN wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.885 0.070 605.955 ;
    END
  END wd_in[164]
  PIN wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.725 0.070 606.795 ;
    END
  END wd_in[165]
  PIN wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.565 0.070 607.635 ;
    END
  END wd_in[166]
  PIN wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.405 0.070 608.475 ;
    END
  END wd_in[167]
  PIN wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.245 0.070 609.315 ;
    END
  END wd_in[168]
  PIN wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.085 0.070 610.155 ;
    END
  END wd_in[169]
  PIN wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.925 0.070 610.995 ;
    END
  END wd_in[170]
  PIN wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.765 0.070 611.835 ;
    END
  END wd_in[171]
  PIN wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.605 0.070 612.675 ;
    END
  END wd_in[172]
  PIN wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.445 0.070 613.515 ;
    END
  END wd_in[173]
  PIN wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.285 0.070 614.355 ;
    END
  END wd_in[174]
  PIN wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.125 0.070 615.195 ;
    END
  END wd_in[175]
  PIN wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.965 0.070 616.035 ;
    END
  END wd_in[176]
  PIN wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.805 0.070 616.875 ;
    END
  END wd_in[177]
  PIN wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.645 0.070 617.715 ;
    END
  END wd_in[178]
  PIN wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.485 0.070 618.555 ;
    END
  END wd_in[179]
  PIN wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.325 0.070 619.395 ;
    END
  END wd_in[180]
  PIN wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.165 0.070 620.235 ;
    END
  END wd_in[181]
  PIN wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.005 0.070 621.075 ;
    END
  END wd_in[182]
  PIN wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.845 0.070 621.915 ;
    END
  END wd_in[183]
  PIN wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.685 0.070 622.755 ;
    END
  END wd_in[184]
  PIN wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.525 0.070 623.595 ;
    END
  END wd_in[185]
  PIN wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.365 0.070 624.435 ;
    END
  END wd_in[186]
  PIN wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.205 0.070 625.275 ;
    END
  END wd_in[187]
  PIN wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.045 0.070 626.115 ;
    END
  END wd_in[188]
  PIN wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.885 0.070 626.955 ;
    END
  END wd_in[189]
  PIN wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.725 0.070 627.795 ;
    END
  END wd_in[190]
  PIN wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.565 0.070 628.635 ;
    END
  END wd_in[191]
  PIN wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.405 0.070 629.475 ;
    END
  END wd_in[192]
  PIN wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.245 0.070 630.315 ;
    END
  END wd_in[193]
  PIN wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.085 0.070 631.155 ;
    END
  END wd_in[194]
  PIN wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.925 0.070 631.995 ;
    END
  END wd_in[195]
  PIN wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.765 0.070 632.835 ;
    END
  END wd_in[196]
  PIN wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.605 0.070 633.675 ;
    END
  END wd_in[197]
  PIN wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.445 0.070 634.515 ;
    END
  END wd_in[198]
  PIN wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.285 0.070 635.355 ;
    END
  END wd_in[199]
  PIN wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.125 0.070 636.195 ;
    END
  END wd_in[200]
  PIN wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.965 0.070 637.035 ;
    END
  END wd_in[201]
  PIN wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.805 0.070 637.875 ;
    END
  END wd_in[202]
  PIN wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.645 0.070 638.715 ;
    END
  END wd_in[203]
  PIN wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.485 0.070 639.555 ;
    END
  END wd_in[204]
  PIN wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.325 0.070 640.395 ;
    END
  END wd_in[205]
  PIN wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.165 0.070 641.235 ;
    END
  END wd_in[206]
  PIN wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.005 0.070 642.075 ;
    END
  END wd_in[207]
  PIN wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.845 0.070 642.915 ;
    END
  END wd_in[208]
  PIN wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.685 0.070 643.755 ;
    END
  END wd_in[209]
  PIN wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.525 0.070 644.595 ;
    END
  END wd_in[210]
  PIN wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.365 0.070 645.435 ;
    END
  END wd_in[211]
  PIN wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.205 0.070 646.275 ;
    END
  END wd_in[212]
  PIN wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.045 0.070 647.115 ;
    END
  END wd_in[213]
  PIN wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.885 0.070 647.955 ;
    END
  END wd_in[214]
  PIN wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.725 0.070 648.795 ;
    END
  END wd_in[215]
  PIN wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.565 0.070 649.635 ;
    END
  END wd_in[216]
  PIN wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.405 0.070 650.475 ;
    END
  END wd_in[217]
  PIN wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.245 0.070 651.315 ;
    END
  END wd_in[218]
  PIN wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.085 0.070 652.155 ;
    END
  END wd_in[219]
  PIN wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.925 0.070 652.995 ;
    END
  END wd_in[220]
  PIN wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.765 0.070 653.835 ;
    END
  END wd_in[221]
  PIN wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.605 0.070 654.675 ;
    END
  END wd_in[222]
  PIN wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.445 0.070 655.515 ;
    END
  END wd_in[223]
  PIN wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.285 0.070 656.355 ;
    END
  END wd_in[224]
  PIN wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.125 0.070 657.195 ;
    END
  END wd_in[225]
  PIN wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.965 0.070 658.035 ;
    END
  END wd_in[226]
  PIN wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.805 0.070 658.875 ;
    END
  END wd_in[227]
  PIN wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.645 0.070 659.715 ;
    END
  END wd_in[228]
  PIN wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.485 0.070 660.555 ;
    END
  END wd_in[229]
  PIN wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.325 0.070 661.395 ;
    END
  END wd_in[230]
  PIN wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.165 0.070 662.235 ;
    END
  END wd_in[231]
  PIN wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.005 0.070 663.075 ;
    END
  END wd_in[232]
  PIN wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.845 0.070 663.915 ;
    END
  END wd_in[233]
  PIN wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.685 0.070 664.755 ;
    END
  END wd_in[234]
  PIN wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.525 0.070 665.595 ;
    END
  END wd_in[235]
  PIN wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.365 0.070 666.435 ;
    END
  END wd_in[236]
  PIN wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.205 0.070 667.275 ;
    END
  END wd_in[237]
  PIN wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.045 0.070 668.115 ;
    END
  END wd_in[238]
  PIN wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.885 0.070 668.955 ;
    END
  END wd_in[239]
  PIN wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.725 0.070 669.795 ;
    END
  END wd_in[240]
  PIN wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.565 0.070 670.635 ;
    END
  END wd_in[241]
  PIN wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.405 0.070 671.475 ;
    END
  END wd_in[242]
  PIN wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.245 0.070 672.315 ;
    END
  END wd_in[243]
  PIN wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.085 0.070 673.155 ;
    END
  END wd_in[244]
  PIN wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.925 0.070 673.995 ;
    END
  END wd_in[245]
  PIN wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.765 0.070 674.835 ;
    END
  END wd_in[246]
  PIN wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.605 0.070 675.675 ;
    END
  END wd_in[247]
  PIN wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.445 0.070 676.515 ;
    END
  END wd_in[248]
  PIN wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.285 0.070 677.355 ;
    END
  END wd_in[249]
  PIN wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.125 0.070 678.195 ;
    END
  END wd_in[250]
  PIN wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.965 0.070 679.035 ;
    END
  END wd_in[251]
  PIN wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.805 0.070 679.875 ;
    END
  END wd_in[252]
  PIN wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.645 0.070 680.715 ;
    END
  END wd_in[253]
  PIN wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.485 0.070 681.555 ;
    END
  END wd_in[254]
  PIN wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.325 0.070 682.395 ;
    END
  END wd_in[255]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.505 0.070 701.575 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.345 0.070 702.415 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.185 0.070 703.255 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.025 0.070 704.095 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.865 0.070 704.935 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.705 0.070 705.775 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.545 0.070 706.615 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.385 0.070 707.455 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.225 0.070 708.295 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.065 0.070 709.135 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.905 0.070 709.975 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.745 0.070 710.815 ;
    END
  END addr_in[11]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.925 0.070 729.995 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.765 0.070 730.835 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.605 0.070 731.675 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 736.400 ;
      RECT 3.500 1.400 3.780 736.400 ;
      RECT 5.740 1.400 6.020 736.400 ;
      RECT 7.980 1.400 8.260 736.400 ;
      RECT 10.220 1.400 10.500 736.400 ;
      RECT 12.460 1.400 12.740 736.400 ;
      RECT 14.700 1.400 14.980 736.400 ;
      RECT 16.940 1.400 17.220 736.400 ;
      RECT 19.180 1.400 19.460 736.400 ;
      RECT 21.420 1.400 21.700 736.400 ;
      RECT 23.660 1.400 23.940 736.400 ;
      RECT 25.900 1.400 26.180 736.400 ;
      RECT 28.140 1.400 28.420 736.400 ;
      RECT 30.380 1.400 30.660 736.400 ;
      RECT 32.620 1.400 32.900 736.400 ;
      RECT 34.860 1.400 35.140 736.400 ;
      RECT 37.100 1.400 37.380 736.400 ;
      RECT 39.340 1.400 39.620 736.400 ;
      RECT 41.580 1.400 41.860 736.400 ;
      RECT 43.820 1.400 44.100 736.400 ;
      RECT 46.060 1.400 46.340 736.400 ;
      RECT 48.300 1.400 48.580 736.400 ;
      RECT 50.540 1.400 50.820 736.400 ;
      RECT 52.780 1.400 53.060 736.400 ;
      RECT 55.020 1.400 55.300 736.400 ;
      RECT 57.260 1.400 57.540 736.400 ;
      RECT 59.500 1.400 59.780 736.400 ;
      RECT 61.740 1.400 62.020 736.400 ;
      RECT 63.980 1.400 64.260 736.400 ;
      RECT 66.220 1.400 66.500 736.400 ;
      RECT 68.460 1.400 68.740 736.400 ;
      RECT 70.700 1.400 70.980 736.400 ;
      RECT 72.940 1.400 73.220 736.400 ;
      RECT 75.180 1.400 75.460 736.400 ;
      RECT 77.420 1.400 77.700 736.400 ;
      RECT 79.660 1.400 79.940 736.400 ;
      RECT 81.900 1.400 82.180 736.400 ;
      RECT 84.140 1.400 84.420 736.400 ;
      RECT 86.380 1.400 86.660 736.400 ;
      RECT 88.620 1.400 88.900 736.400 ;
      RECT 90.860 1.400 91.140 736.400 ;
      RECT 93.100 1.400 93.380 736.400 ;
      RECT 95.340 1.400 95.620 736.400 ;
      RECT 97.580 1.400 97.860 736.400 ;
      RECT 99.820 1.400 100.100 736.400 ;
      RECT 102.060 1.400 102.340 736.400 ;
      RECT 104.300 1.400 104.580 736.400 ;
      RECT 106.540 1.400 106.820 736.400 ;
      RECT 108.780 1.400 109.060 736.400 ;
      RECT 111.020 1.400 111.300 736.400 ;
      RECT 113.260 1.400 113.540 736.400 ;
      RECT 115.500 1.400 115.780 736.400 ;
      RECT 117.740 1.400 118.020 736.400 ;
      RECT 119.980 1.400 120.260 736.400 ;
      RECT 122.220 1.400 122.500 736.400 ;
      RECT 124.460 1.400 124.740 736.400 ;
      RECT 126.700 1.400 126.980 736.400 ;
      RECT 128.940 1.400 129.220 736.400 ;
      RECT 131.180 1.400 131.460 736.400 ;
      RECT 133.420 1.400 133.700 736.400 ;
      RECT 135.660 1.400 135.940 736.400 ;
      RECT 137.900 1.400 138.180 736.400 ;
      RECT 140.140 1.400 140.420 736.400 ;
      RECT 142.380 1.400 142.660 736.400 ;
      RECT 144.620 1.400 144.900 736.400 ;
      RECT 146.860 1.400 147.140 736.400 ;
      RECT 149.100 1.400 149.380 736.400 ;
      RECT 151.340 1.400 151.620 736.400 ;
      RECT 153.580 1.400 153.860 736.400 ;
      RECT 155.820 1.400 156.100 736.400 ;
      RECT 158.060 1.400 158.340 736.400 ;
      RECT 160.300 1.400 160.580 736.400 ;
      RECT 162.540 1.400 162.820 736.400 ;
      RECT 164.780 1.400 165.060 736.400 ;
      RECT 167.020 1.400 167.300 736.400 ;
      RECT 169.260 1.400 169.540 736.400 ;
      RECT 171.500 1.400 171.780 736.400 ;
      RECT 173.740 1.400 174.020 736.400 ;
      RECT 175.980 1.400 176.260 736.400 ;
      RECT 178.220 1.400 178.500 736.400 ;
      RECT 180.460 1.400 180.740 736.400 ;
      RECT 182.700 1.400 182.980 736.400 ;
      RECT 184.940 1.400 185.220 736.400 ;
      RECT 187.180 1.400 187.460 736.400 ;
      RECT 189.420 1.400 189.700 736.400 ;
      RECT 191.660 1.400 191.940 736.400 ;
      RECT 193.900 1.400 194.180 736.400 ;
      RECT 196.140 1.400 196.420 736.400 ;
      RECT 198.380 1.400 198.660 736.400 ;
      RECT 200.620 1.400 200.900 736.400 ;
      RECT 202.860 1.400 203.140 736.400 ;
      RECT 205.100 1.400 205.380 736.400 ;
      RECT 207.340 1.400 207.620 736.400 ;
      RECT 209.580 1.400 209.860 736.400 ;
      RECT 211.820 1.400 212.100 736.400 ;
      RECT 214.060 1.400 214.340 736.400 ;
      RECT 216.300 1.400 216.580 736.400 ;
      RECT 218.540 1.400 218.820 736.400 ;
      RECT 220.780 1.400 221.060 736.400 ;
      RECT 223.020 1.400 223.300 736.400 ;
      RECT 225.260 1.400 225.540 736.400 ;
      RECT 227.500 1.400 227.780 736.400 ;
      RECT 229.740 1.400 230.020 736.400 ;
      RECT 231.980 1.400 232.260 736.400 ;
      RECT 234.220 1.400 234.500 736.400 ;
      RECT 236.460 1.400 236.740 736.400 ;
      RECT 238.700 1.400 238.980 736.400 ;
      RECT 240.940 1.400 241.220 736.400 ;
      RECT 243.180 1.400 243.460 736.400 ;
      RECT 245.420 1.400 245.700 736.400 ;
      RECT 247.660 1.400 247.940 736.400 ;
      RECT 249.900 1.400 250.180 736.400 ;
      RECT 252.140 1.400 252.420 736.400 ;
      RECT 254.380 1.400 254.660 736.400 ;
      RECT 256.620 1.400 256.900 736.400 ;
      RECT 258.860 1.400 259.140 736.400 ;
      RECT 261.100 1.400 261.380 736.400 ;
      RECT 263.340 1.400 263.620 736.400 ;
      RECT 265.580 1.400 265.860 736.400 ;
      RECT 267.820 1.400 268.100 736.400 ;
      RECT 270.060 1.400 270.340 736.400 ;
      RECT 272.300 1.400 272.580 736.400 ;
      RECT 274.540 1.400 274.820 736.400 ;
      RECT 276.780 1.400 277.060 736.400 ;
      RECT 279.020 1.400 279.300 736.400 ;
      RECT 281.260 1.400 281.540 736.400 ;
      RECT 283.500 1.400 283.780 736.400 ;
      RECT 285.740 1.400 286.020 736.400 ;
      RECT 287.980 1.400 288.260 736.400 ;
      RECT 290.220 1.400 290.500 736.400 ;
      RECT 292.460 1.400 292.740 736.400 ;
      RECT 294.700 1.400 294.980 736.400 ;
      RECT 296.940 1.400 297.220 736.400 ;
      RECT 299.180 1.400 299.460 736.400 ;
      RECT 301.420 1.400 301.700 736.400 ;
      RECT 303.660 1.400 303.940 736.400 ;
      RECT 305.900 1.400 306.180 736.400 ;
      RECT 308.140 1.400 308.420 736.400 ;
      RECT 310.380 1.400 310.660 736.400 ;
      RECT 312.620 1.400 312.900 736.400 ;
      RECT 314.860 1.400 315.140 736.400 ;
      RECT 317.100 1.400 317.380 736.400 ;
      RECT 319.340 1.400 319.620 736.400 ;
      RECT 321.580 1.400 321.860 736.400 ;
      RECT 323.820 1.400 324.100 736.400 ;
      RECT 326.060 1.400 326.340 736.400 ;
      RECT 328.300 1.400 328.580 736.400 ;
      RECT 330.540 1.400 330.820 736.400 ;
      RECT 332.780 1.400 333.060 736.400 ;
      RECT 335.020 1.400 335.300 736.400 ;
      RECT 337.260 1.400 337.540 736.400 ;
      RECT 339.500 1.400 339.780 736.400 ;
      RECT 341.740 1.400 342.020 736.400 ;
      RECT 343.980 1.400 344.260 736.400 ;
      RECT 346.220 1.400 346.500 736.400 ;
      RECT 348.460 1.400 348.740 736.400 ;
      RECT 350.700 1.400 350.980 736.400 ;
      RECT 352.940 1.400 353.220 736.400 ;
      RECT 355.180 1.400 355.460 736.400 ;
      RECT 357.420 1.400 357.700 736.400 ;
      RECT 359.660 1.400 359.940 736.400 ;
      RECT 361.900 1.400 362.180 736.400 ;
      RECT 364.140 1.400 364.420 736.400 ;
      RECT 366.380 1.400 366.660 736.400 ;
      RECT 368.620 1.400 368.900 736.400 ;
      RECT 370.860 1.400 371.140 736.400 ;
      RECT 373.100 1.400 373.380 736.400 ;
      RECT 375.340 1.400 375.620 736.400 ;
      RECT 377.580 1.400 377.860 736.400 ;
      RECT 379.820 1.400 380.100 736.400 ;
      RECT 382.060 1.400 382.340 736.400 ;
      RECT 384.300 1.400 384.580 736.400 ;
      RECT 386.540 1.400 386.820 736.400 ;
      RECT 388.780 1.400 389.060 736.400 ;
      RECT 391.020 1.400 391.300 736.400 ;
      RECT 393.260 1.400 393.540 736.400 ;
      RECT 395.500 1.400 395.780 736.400 ;
      RECT 397.740 1.400 398.020 736.400 ;
      RECT 399.980 1.400 400.260 736.400 ;
      RECT 402.220 1.400 402.500 736.400 ;
      RECT 404.460 1.400 404.740 736.400 ;
      RECT 406.700 1.400 406.980 736.400 ;
      RECT 408.940 1.400 409.220 736.400 ;
      RECT 411.180 1.400 411.460 736.400 ;
      RECT 413.420 1.400 413.700 736.400 ;
      RECT 415.660 1.400 415.940 736.400 ;
      RECT 417.900 1.400 418.180 736.400 ;
      RECT 420.140 1.400 420.420 736.400 ;
      RECT 422.380 1.400 422.660 736.400 ;
      RECT 424.620 1.400 424.900 736.400 ;
      RECT 426.860 1.400 427.140 736.400 ;
      RECT 429.100 1.400 429.380 736.400 ;
      RECT 431.340 1.400 431.620 736.400 ;
      RECT 433.580 1.400 433.860 736.400 ;
      RECT 435.820 1.400 436.100 736.400 ;
      RECT 438.060 1.400 438.340 736.400 ;
      RECT 440.300 1.400 440.580 736.400 ;
      RECT 442.540 1.400 442.820 736.400 ;
      RECT 444.780 1.400 445.060 736.400 ;
      RECT 447.020 1.400 447.300 736.400 ;
      RECT 449.260 1.400 449.540 736.400 ;
      RECT 451.500 1.400 451.780 736.400 ;
      RECT 453.740 1.400 454.020 736.400 ;
      RECT 455.980 1.400 456.260 736.400 ;
      RECT 458.220 1.400 458.500 736.400 ;
      RECT 460.460 1.400 460.740 736.400 ;
      RECT 462.700 1.400 462.980 736.400 ;
      RECT 464.940 1.400 465.220 736.400 ;
      RECT 467.180 1.400 467.460 736.400 ;
      RECT 469.420 1.400 469.700 736.400 ;
      RECT 471.660 1.400 471.940 736.400 ;
      RECT 473.900 1.400 474.180 736.400 ;
      RECT 476.140 1.400 476.420 736.400 ;
      RECT 478.380 1.400 478.660 736.400 ;
      RECT 480.620 1.400 480.900 736.400 ;
      RECT 482.860 1.400 483.140 736.400 ;
      RECT 485.100 1.400 485.380 736.400 ;
      RECT 487.340 1.400 487.620 736.400 ;
      RECT 489.580 1.400 489.860 736.400 ;
      RECT 491.820 1.400 492.100 736.400 ;
      RECT 494.060 1.400 494.340 736.400 ;
      RECT 496.300 1.400 496.580 736.400 ;
      RECT 498.540 1.400 498.820 736.400 ;
      RECT 500.780 1.400 501.060 736.400 ;
      RECT 503.020 1.400 503.300 736.400 ;
      RECT 505.260 1.400 505.540 736.400 ;
      RECT 507.500 1.400 507.780 736.400 ;
      RECT 509.740 1.400 510.020 736.400 ;
      RECT 511.980 1.400 512.260 736.400 ;
      RECT 514.220 1.400 514.500 736.400 ;
      RECT 516.460 1.400 516.740 736.400 ;
      RECT 518.700 1.400 518.980 736.400 ;
      RECT 520.940 1.400 521.220 736.400 ;
      RECT 523.180 1.400 523.460 736.400 ;
      RECT 525.420 1.400 525.700 736.400 ;
      RECT 527.660 1.400 527.940 736.400 ;
      RECT 529.900 1.400 530.180 736.400 ;
      RECT 532.140 1.400 532.420 736.400 ;
      RECT 534.380 1.400 534.660 736.400 ;
      RECT 536.620 1.400 536.900 736.400 ;
      RECT 538.860 1.400 539.140 736.400 ;
      RECT 541.100 1.400 541.380 736.400 ;
      RECT 543.340 1.400 543.620 736.400 ;
      RECT 545.580 1.400 545.860 736.400 ;
      RECT 547.820 1.400 548.100 736.400 ;
      RECT 550.060 1.400 550.340 736.400 ;
      RECT 552.300 1.400 552.580 736.400 ;
      RECT 554.540 1.400 554.820 736.400 ;
      RECT 556.780 1.400 557.060 736.400 ;
      RECT 559.020 1.400 559.300 736.400 ;
      RECT 561.260 1.400 561.540 736.400 ;
      RECT 563.500 1.400 563.780 736.400 ;
      RECT 565.740 1.400 566.020 736.400 ;
      RECT 567.980 1.400 568.260 736.400 ;
      RECT 570.220 1.400 570.500 736.400 ;
      RECT 572.460 1.400 572.740 736.400 ;
      RECT 574.700 1.400 574.980 736.400 ;
      RECT 576.940 1.400 577.220 736.400 ;
      RECT 579.180 1.400 579.460 736.400 ;
      RECT 581.420 1.400 581.700 736.400 ;
      RECT 583.660 1.400 583.940 736.400 ;
      RECT 585.900 1.400 586.180 736.400 ;
      RECT 588.140 1.400 588.420 736.400 ;
      RECT 590.380 1.400 590.660 736.400 ;
      RECT 592.620 1.400 592.900 736.400 ;
      RECT 594.860 1.400 595.140 736.400 ;
      RECT 597.100 1.400 597.380 736.400 ;
      RECT 599.340 1.400 599.620 736.400 ;
      RECT 601.580 1.400 601.860 736.400 ;
      RECT 603.820 1.400 604.100 736.400 ;
      RECT 606.060 1.400 606.340 736.400 ;
      RECT 608.300 1.400 608.580 736.400 ;
      RECT 610.540 1.400 610.820 736.400 ;
      RECT 612.780 1.400 613.060 736.400 ;
      RECT 615.020 1.400 615.300 736.400 ;
      RECT 617.260 1.400 617.540 736.400 ;
      RECT 619.500 1.400 619.780 736.400 ;
      RECT 621.740 1.400 622.020 736.400 ;
      RECT 623.980 1.400 624.260 736.400 ;
      RECT 626.220 1.400 626.500 736.400 ;
      RECT 628.460 1.400 628.740 736.400 ;
      RECT 630.700 1.400 630.980 736.400 ;
      RECT 632.940 1.400 633.220 736.400 ;
      RECT 635.180 1.400 635.460 736.400 ;
      RECT 637.420 1.400 637.700 736.400 ;
      RECT 639.660 1.400 639.940 736.400 ;
      RECT 641.900 1.400 642.180 736.400 ;
      RECT 644.140 1.400 644.420 736.400 ;
      RECT 646.380 1.400 646.660 736.400 ;
      RECT 648.620 1.400 648.900 736.400 ;
      RECT 650.860 1.400 651.140 736.400 ;
      RECT 653.100 1.400 653.380 736.400 ;
      RECT 655.340 1.400 655.620 736.400 ;
      RECT 657.580 1.400 657.860 736.400 ;
      RECT 659.820 1.400 660.100 736.400 ;
      RECT 662.060 1.400 662.340 736.400 ;
      RECT 664.300 1.400 664.580 736.400 ;
      RECT 666.540 1.400 666.820 736.400 ;
      RECT 668.780 1.400 669.060 736.400 ;
      RECT 671.020 1.400 671.300 736.400 ;
      RECT 673.260 1.400 673.540 736.400 ;
      RECT 675.500 1.400 675.780 736.400 ;
      RECT 677.740 1.400 678.020 736.400 ;
      RECT 679.980 1.400 680.260 736.400 ;
      RECT 682.220 1.400 682.500 736.400 ;
      RECT 684.460 1.400 684.740 736.400 ;
      RECT 686.700 1.400 686.980 736.400 ;
      RECT 688.940 1.400 689.220 736.400 ;
      RECT 691.180 1.400 691.460 736.400 ;
      RECT 693.420 1.400 693.700 736.400 ;
      RECT 695.660 1.400 695.940 736.400 ;
      RECT 697.900 1.400 698.180 736.400 ;
      RECT 700.140 1.400 700.420 736.400 ;
      RECT 702.380 1.400 702.660 736.400 ;
      RECT 704.620 1.400 704.900 736.400 ;
      RECT 706.860 1.400 707.140 736.400 ;
      RECT 709.100 1.400 709.380 736.400 ;
      RECT 711.340 1.400 711.620 736.400 ;
      RECT 713.580 1.400 713.860 736.400 ;
      RECT 715.820 1.400 716.100 736.400 ;
      RECT 718.060 1.400 718.340 736.400 ;
      RECT 720.300 1.400 720.580 736.400 ;
      RECT 722.540 1.400 722.820 736.400 ;
      RECT 724.780 1.400 725.060 736.400 ;
      RECT 727.020 1.400 727.300 736.400 ;
      RECT 729.260 1.400 729.540 736.400 ;
      RECT 731.500 1.400 731.780 736.400 ;
      RECT 733.740 1.400 734.020 736.400 ;
      RECT 735.980 1.400 736.260 736.400 ;
      RECT 738.220 1.400 738.500 736.400 ;
      RECT 740.460 1.400 740.740 736.400 ;
      RECT 742.700 1.400 742.980 736.400 ;
      RECT 744.940 1.400 745.220 736.400 ;
      RECT 747.180 1.400 747.460 736.400 ;
      RECT 749.420 1.400 749.700 736.400 ;
      RECT 751.660 1.400 751.940 736.400 ;
      RECT 753.900 1.400 754.180 736.400 ;
      RECT 756.140 1.400 756.420 736.400 ;
      RECT 758.380 1.400 758.660 736.400 ;
      RECT 760.620 1.400 760.900 736.400 ;
      RECT 762.860 1.400 763.140 736.400 ;
      RECT 765.100 1.400 765.380 736.400 ;
      RECT 767.340 1.400 767.620 736.400 ;
      RECT 769.580 1.400 769.860 736.400 ;
      RECT 771.820 1.400 772.100 736.400 ;
      RECT 774.060 1.400 774.340 736.400 ;
      RECT 776.300 1.400 776.580 736.400 ;
      RECT 778.540 1.400 778.820 736.400 ;
      RECT 780.780 1.400 781.060 736.400 ;
      RECT 783.020 1.400 783.300 736.400 ;
      RECT 785.260 1.400 785.540 736.400 ;
      RECT 787.500 1.400 787.780 736.400 ;
      RECT 789.740 1.400 790.020 736.400 ;
      RECT 791.980 1.400 792.260 736.400 ;
      RECT 794.220 1.400 794.500 736.400 ;
      RECT 796.460 1.400 796.740 736.400 ;
      RECT 798.700 1.400 798.980 736.400 ;
      RECT 800.940 1.400 801.220 736.400 ;
      RECT 803.180 1.400 803.460 736.400 ;
      RECT 805.420 1.400 805.700 736.400 ;
      RECT 807.660 1.400 807.940 736.400 ;
      RECT 809.900 1.400 810.180 736.400 ;
      RECT 812.140 1.400 812.420 736.400 ;
      RECT 814.380 1.400 814.660 736.400 ;
      RECT 816.620 1.400 816.900 736.400 ;
      RECT 818.860 1.400 819.140 736.400 ;
      RECT 821.100 1.400 821.380 736.400 ;
      RECT 823.340 1.400 823.620 736.400 ;
      RECT 825.580 1.400 825.860 736.400 ;
      RECT 827.820 1.400 828.100 736.400 ;
      RECT 830.060 1.400 830.340 736.400 ;
      RECT 832.300 1.400 832.580 736.400 ;
      RECT 834.540 1.400 834.820 736.400 ;
      RECT 836.780 1.400 837.060 736.400 ;
      RECT 839.020 1.400 839.300 736.400 ;
      RECT 841.260 1.400 841.540 736.400 ;
      RECT 843.500 1.400 843.780 736.400 ;
      RECT 845.740 1.400 846.020 736.400 ;
      RECT 847.980 1.400 848.260 736.400 ;
      RECT 850.220 1.400 850.500 736.400 ;
      RECT 852.460 1.400 852.740 736.400 ;
      RECT 854.700 1.400 854.980 736.400 ;
      RECT 856.940 1.400 857.220 736.400 ;
      RECT 859.180 1.400 859.460 736.400 ;
      RECT 861.420 1.400 861.700 736.400 ;
      RECT 863.660 1.400 863.940 736.400 ;
      RECT 865.900 1.400 866.180 736.400 ;
      RECT 868.140 1.400 868.420 736.400 ;
      RECT 870.380 1.400 870.660 736.400 ;
      RECT 872.620 1.400 872.900 736.400 ;
      RECT 874.860 1.400 875.140 736.400 ;
      RECT 877.100 1.400 877.380 736.400 ;
      RECT 879.340 1.400 879.620 736.400 ;
      RECT 881.580 1.400 881.860 736.400 ;
      RECT 883.820 1.400 884.100 736.400 ;
      RECT 886.060 1.400 886.340 736.400 ;
      RECT 888.300 1.400 888.580 736.400 ;
      RECT 890.540 1.400 890.820 736.400 ;
      RECT 892.780 1.400 893.060 736.400 ;
      RECT 895.020 1.400 895.300 736.400 ;
      RECT 897.260 1.400 897.540 736.400 ;
      RECT 899.500 1.400 899.780 736.400 ;
      RECT 901.740 1.400 902.020 736.400 ;
      RECT 903.980 1.400 904.260 736.400 ;
      RECT 906.220 1.400 906.500 736.400 ;
      RECT 908.460 1.400 908.740 736.400 ;
      RECT 910.700 1.400 910.980 736.400 ;
      RECT 912.940 1.400 913.220 736.400 ;
      RECT 915.180 1.400 915.460 736.400 ;
      RECT 917.420 1.400 917.700 736.400 ;
      RECT 919.660 1.400 919.940 736.400 ;
      RECT 921.900 1.400 922.180 736.400 ;
      RECT 924.140 1.400 924.420 736.400 ;
      RECT 926.380 1.400 926.660 736.400 ;
      RECT 928.620 1.400 928.900 736.400 ;
      RECT 930.860 1.400 931.140 736.400 ;
      RECT 933.100 1.400 933.380 736.400 ;
      RECT 935.340 1.400 935.620 736.400 ;
      RECT 937.580 1.400 937.860 736.400 ;
      RECT 939.820 1.400 940.100 736.400 ;
      RECT 942.060 1.400 942.340 736.400 ;
      RECT 944.300 1.400 944.580 736.400 ;
      RECT 946.540 1.400 946.820 736.400 ;
      RECT 948.780 1.400 949.060 736.400 ;
      RECT 951.020 1.400 951.300 736.400 ;
      RECT 953.260 1.400 953.540 736.400 ;
      RECT 955.500 1.400 955.780 736.400 ;
      RECT 957.740 1.400 958.020 736.400 ;
      RECT 959.980 1.400 960.260 736.400 ;
      RECT 962.220 1.400 962.500 736.400 ;
      RECT 964.460 1.400 964.740 736.400 ;
      RECT 966.700 1.400 966.980 736.400 ;
      RECT 968.940 1.400 969.220 736.400 ;
      RECT 971.180 1.400 971.460 736.400 ;
      RECT 973.420 1.400 973.700 736.400 ;
      RECT 975.660 1.400 975.940 736.400 ;
      RECT 977.900 1.400 978.180 736.400 ;
      RECT 980.140 1.400 980.420 736.400 ;
      RECT 982.380 1.400 982.660 736.400 ;
      RECT 984.620 1.400 984.900 736.400 ;
      RECT 986.860 1.400 987.140 736.400 ;
      RECT 989.100 1.400 989.380 736.400 ;
      RECT 991.340 1.400 991.620 736.400 ;
      RECT 993.580 1.400 993.860 736.400 ;
      RECT 995.820 1.400 996.100 736.400 ;
      RECT 998.060 1.400 998.340 736.400 ;
      RECT 1000.300 1.400 1000.580 736.400 ;
      RECT 1002.540 1.400 1002.820 736.400 ;
      RECT 1004.780 1.400 1005.060 736.400 ;
      RECT 1007.020 1.400 1007.300 736.400 ;
      RECT 1009.260 1.400 1009.540 736.400 ;
      RECT 1011.500 1.400 1011.780 736.400 ;
      RECT 1013.740 1.400 1014.020 736.400 ;
      RECT 1015.980 1.400 1016.260 736.400 ;
      RECT 1018.220 1.400 1018.500 736.400 ;
      RECT 1020.460 1.400 1020.740 736.400 ;
      RECT 1022.700 1.400 1022.980 736.400 ;
      RECT 1024.940 1.400 1025.220 736.400 ;
      RECT 1027.180 1.400 1027.460 736.400 ;
      RECT 1029.420 1.400 1029.700 736.400 ;
      RECT 1031.660 1.400 1031.940 736.400 ;
      RECT 1033.900 1.400 1034.180 736.400 ;
      RECT 1036.140 1.400 1036.420 736.400 ;
      RECT 1038.380 1.400 1038.660 736.400 ;
      RECT 1040.620 1.400 1040.900 736.400 ;
      RECT 1042.860 1.400 1043.140 736.400 ;
      RECT 1045.100 1.400 1045.380 736.400 ;
      RECT 1047.340 1.400 1047.620 736.400 ;
      RECT 1049.580 1.400 1049.860 736.400 ;
      RECT 1051.820 1.400 1052.100 736.400 ;
      RECT 1054.060 1.400 1054.340 736.400 ;
      RECT 1056.300 1.400 1056.580 736.400 ;
      RECT 1058.540 1.400 1058.820 736.400 ;
      RECT 1060.780 1.400 1061.060 736.400 ;
      RECT 1063.020 1.400 1063.300 736.400 ;
      RECT 1065.260 1.400 1065.540 736.400 ;
      RECT 1067.500 1.400 1067.780 736.400 ;
      RECT 1069.740 1.400 1070.020 736.400 ;
      RECT 1071.980 1.400 1072.260 736.400 ;
      RECT 1074.220 1.400 1074.500 736.400 ;
      RECT 1076.460 1.400 1076.740 736.400 ;
      RECT 1078.700 1.400 1078.980 736.400 ;
      RECT 1080.940 1.400 1081.220 736.400 ;
      RECT 1083.180 1.400 1083.460 736.400 ;
      RECT 1085.420 1.400 1085.700 736.400 ;
      RECT 1087.660 1.400 1087.940 736.400 ;
      RECT 1089.900 1.400 1090.180 736.400 ;
      RECT 1092.140 1.400 1092.420 736.400 ;
      RECT 1094.380 1.400 1094.660 736.400 ;
      RECT 1096.620 1.400 1096.900 736.400 ;
      RECT 1098.860 1.400 1099.140 736.400 ;
      RECT 1101.100 1.400 1101.380 736.400 ;
      RECT 1103.340 1.400 1103.620 736.400 ;
      RECT 1105.580 1.400 1105.860 736.400 ;
      RECT 1107.820 1.400 1108.100 736.400 ;
      RECT 1110.060 1.400 1110.340 736.400 ;
      RECT 1112.300 1.400 1112.580 736.400 ;
      RECT 1114.540 1.400 1114.820 736.400 ;
      RECT 1116.780 1.400 1117.060 736.400 ;
      RECT 1119.020 1.400 1119.300 736.400 ;
      RECT 1121.260 1.400 1121.540 736.400 ;
      RECT 1123.500 1.400 1123.780 736.400 ;
      RECT 1125.740 1.400 1126.020 736.400 ;
      RECT 1127.980 1.400 1128.260 736.400 ;
      RECT 1130.220 1.400 1130.500 736.400 ;
      RECT 1132.460 1.400 1132.740 736.400 ;
      RECT 1134.700 1.400 1134.980 736.400 ;
      RECT 1136.940 1.400 1137.220 736.400 ;
      RECT 1139.180 1.400 1139.460 736.400 ;
      RECT 1141.420 1.400 1141.700 736.400 ;
      RECT 1143.660 1.400 1143.940 736.400 ;
      RECT 1145.900 1.400 1146.180 736.400 ;
      RECT 1148.140 1.400 1148.420 736.400 ;
      RECT 1150.380 1.400 1150.660 736.400 ;
      RECT 1152.620 1.400 1152.900 736.400 ;
      RECT 1154.860 1.400 1155.140 736.400 ;
      RECT 1157.100 1.400 1157.380 736.400 ;
      RECT 1159.340 1.400 1159.620 736.400 ;
      RECT 1161.580 1.400 1161.860 736.400 ;
      RECT 1163.820 1.400 1164.100 736.400 ;
      RECT 1166.060 1.400 1166.340 736.400 ;
      RECT 1168.300 1.400 1168.580 736.400 ;
      RECT 1170.540 1.400 1170.820 736.400 ;
      RECT 1172.780 1.400 1173.060 736.400 ;
      RECT 1175.020 1.400 1175.300 736.400 ;
      RECT 1177.260 1.400 1177.540 736.400 ;
      RECT 1179.500 1.400 1179.780 736.400 ;
      RECT 1181.740 1.400 1182.020 736.400 ;
      RECT 1183.980 1.400 1184.260 736.400 ;
      RECT 1186.220 1.400 1186.500 736.400 ;
      RECT 1188.460 1.400 1188.740 736.400 ;
      RECT 1190.700 1.400 1190.980 736.400 ;
      RECT 1192.940 1.400 1193.220 736.400 ;
      RECT 1195.180 1.400 1195.460 736.400 ;
      RECT 1197.420 1.400 1197.700 736.400 ;
      RECT 1199.660 1.400 1199.940 736.400 ;
      RECT 1201.900 1.400 1202.180 736.400 ;
      RECT 1204.140 1.400 1204.420 736.400 ;
      RECT 1206.380 1.400 1206.660 736.400 ;
      RECT 1208.620 1.400 1208.900 736.400 ;
      RECT 1210.860 1.400 1211.140 736.400 ;
      RECT 1213.100 1.400 1213.380 736.400 ;
      RECT 1215.340 1.400 1215.620 736.400 ;
      RECT 1217.580 1.400 1217.860 736.400 ;
      RECT 1219.820 1.400 1220.100 736.400 ;
      RECT 1222.060 1.400 1222.340 736.400 ;
      RECT 1224.300 1.400 1224.580 736.400 ;
      RECT 1226.540 1.400 1226.820 736.400 ;
      RECT 1228.780 1.400 1229.060 736.400 ;
      RECT 1231.020 1.400 1231.300 736.400 ;
      RECT 1233.260 1.400 1233.540 736.400 ;
      RECT 1235.500 1.400 1235.780 736.400 ;
      RECT 1237.740 1.400 1238.020 736.400 ;
      RECT 1239.980 1.400 1240.260 736.400 ;
      RECT 1242.220 1.400 1242.500 736.400 ;
      RECT 1244.460 1.400 1244.740 736.400 ;
      RECT 1246.700 1.400 1246.980 736.400 ;
      RECT 1248.940 1.400 1249.220 736.400 ;
      RECT 1251.180 1.400 1251.460 736.400 ;
      RECT 1253.420 1.400 1253.700 736.400 ;
      RECT 1255.660 1.400 1255.940 736.400 ;
      RECT 1257.900 1.400 1258.180 736.400 ;
      RECT 1260.140 1.400 1260.420 736.400 ;
      RECT 1262.380 1.400 1262.660 736.400 ;
      RECT 1264.620 1.400 1264.900 736.400 ;
      RECT 1266.860 1.400 1267.140 736.400 ;
      RECT 1269.100 1.400 1269.380 736.400 ;
      RECT 1271.340 1.400 1271.620 736.400 ;
      RECT 1273.580 1.400 1273.860 736.400 ;
      RECT 1275.820 1.400 1276.100 736.400 ;
      RECT 1278.060 1.400 1278.340 736.400 ;
      RECT 1280.300 1.400 1280.580 736.400 ;
      RECT 1282.540 1.400 1282.820 736.400 ;
      RECT 1284.780 1.400 1285.060 736.400 ;
      RECT 1287.020 1.400 1287.300 736.400 ;
      RECT 1289.260 1.400 1289.540 736.400 ;
      RECT 1291.500 1.400 1291.780 736.400 ;
      RECT 1293.740 1.400 1294.020 736.400 ;
      RECT 1295.980 1.400 1296.260 736.400 ;
      RECT 1298.220 1.400 1298.500 736.400 ;
      RECT 1300.460 1.400 1300.740 736.400 ;
      RECT 1302.700 1.400 1302.980 736.400 ;
      RECT 1304.940 1.400 1305.220 736.400 ;
      RECT 1307.180 1.400 1307.460 736.400 ;
      RECT 1309.420 1.400 1309.700 736.400 ;
      RECT 1311.660 1.400 1311.940 736.400 ;
      RECT 1313.900 1.400 1314.180 736.400 ;
      RECT 1316.140 1.400 1316.420 736.400 ;
      RECT 1318.380 1.400 1318.660 736.400 ;
      RECT 1320.620 1.400 1320.900 736.400 ;
      RECT 1322.860 1.400 1323.140 736.400 ;
      RECT 1325.100 1.400 1325.380 736.400 ;
      RECT 1327.340 1.400 1327.620 736.400 ;
      RECT 1329.580 1.400 1329.860 736.400 ;
      RECT 1331.820 1.400 1332.100 736.400 ;
      RECT 1334.060 1.400 1334.340 736.400 ;
      RECT 1336.300 1.400 1336.580 736.400 ;
      RECT 1338.540 1.400 1338.820 736.400 ;
      RECT 1340.780 1.400 1341.060 736.400 ;
      RECT 1343.020 1.400 1343.300 736.400 ;
      RECT 1345.260 1.400 1345.540 736.400 ;
      RECT 1347.500 1.400 1347.780 736.400 ;
      RECT 1349.740 1.400 1350.020 736.400 ;
      RECT 1351.980 1.400 1352.260 736.400 ;
      RECT 1354.220 1.400 1354.500 736.400 ;
      RECT 1356.460 1.400 1356.740 736.400 ;
      RECT 1358.700 1.400 1358.980 736.400 ;
      RECT 1360.940 1.400 1361.220 736.400 ;
      RECT 1363.180 1.400 1363.460 736.400 ;
      RECT 1365.420 1.400 1365.700 736.400 ;
      RECT 1367.660 1.400 1367.940 736.400 ;
      RECT 1369.900 1.400 1370.180 736.400 ;
      RECT 1372.140 1.400 1372.420 736.400 ;
      RECT 1374.380 1.400 1374.660 736.400 ;
      RECT 1376.620 1.400 1376.900 736.400 ;
      RECT 1378.860 1.400 1379.140 736.400 ;
      RECT 1381.100 1.400 1381.380 736.400 ;
      RECT 1383.340 1.400 1383.620 736.400 ;
      RECT 1385.580 1.400 1385.860 736.400 ;
      RECT 1387.820 1.400 1388.100 736.400 ;
      RECT 1390.060 1.400 1390.340 736.400 ;
      RECT 1392.300 1.400 1392.580 736.400 ;
      RECT 1394.540 1.400 1394.820 736.400 ;
      RECT 1396.780 1.400 1397.060 736.400 ;
      RECT 1399.020 1.400 1399.300 736.400 ;
      RECT 1401.260 1.400 1401.540 736.400 ;
      RECT 1403.500 1.400 1403.780 736.400 ;
      RECT 1405.740 1.400 1406.020 736.400 ;
      RECT 1407.980 1.400 1408.260 736.400 ;
      RECT 1410.220 1.400 1410.500 736.400 ;
      RECT 1412.460 1.400 1412.740 736.400 ;
      RECT 1414.700 1.400 1414.980 736.400 ;
      RECT 1416.940 1.400 1417.220 736.400 ;
      RECT 1419.180 1.400 1419.460 736.400 ;
      RECT 1421.420 1.400 1421.700 736.400 ;
      RECT 1423.660 1.400 1423.940 736.400 ;
      RECT 1425.900 1.400 1426.180 736.400 ;
      RECT 1428.140 1.400 1428.420 736.400 ;
      RECT 1430.380 1.400 1430.660 736.400 ;
      RECT 1432.620 1.400 1432.900 736.400 ;
      RECT 1434.860 1.400 1435.140 736.400 ;
      RECT 1437.100 1.400 1437.380 736.400 ;
      RECT 1439.340 1.400 1439.620 736.400 ;
      RECT 1441.580 1.400 1441.860 736.400 ;
      RECT 1443.820 1.400 1444.100 736.400 ;
      RECT 1446.060 1.400 1446.340 736.400 ;
      RECT 1448.300 1.400 1448.580 736.400 ;
      RECT 1450.540 1.400 1450.820 736.400 ;
      RECT 1452.780 1.400 1453.060 736.400 ;
      RECT 1455.020 1.400 1455.300 736.400 ;
      RECT 1457.260 1.400 1457.540 736.400 ;
      RECT 1459.500 1.400 1459.780 736.400 ;
      RECT 1461.740 1.400 1462.020 736.400 ;
      RECT 1463.980 1.400 1464.260 736.400 ;
      RECT 1466.220 1.400 1466.500 736.400 ;
      RECT 1468.460 1.400 1468.740 736.400 ;
      RECT 1470.700 1.400 1470.980 736.400 ;
      RECT 1472.940 1.400 1473.220 736.400 ;
      RECT 1475.180 1.400 1475.460 736.400 ;
      RECT 1477.420 1.400 1477.700 736.400 ;
      RECT 1479.660 1.400 1479.940 736.400 ;
      RECT 1481.900 1.400 1482.180 736.400 ;
      RECT 1484.140 1.400 1484.420 736.400 ;
      RECT 1486.380 1.400 1486.660 736.400 ;
      RECT 1488.620 1.400 1488.900 736.400 ;
      RECT 1490.860 1.400 1491.140 736.400 ;
      RECT 1493.100 1.400 1493.380 736.400 ;
      RECT 1495.340 1.400 1495.620 736.400 ;
      RECT 1497.580 1.400 1497.860 736.400 ;
      RECT 1499.820 1.400 1500.100 736.400 ;
      RECT 1502.060 1.400 1502.340 736.400 ;
      RECT 1504.300 1.400 1504.580 736.400 ;
      RECT 1506.540 1.400 1506.820 736.400 ;
      RECT 1508.780 1.400 1509.060 736.400 ;
      RECT 1511.020 1.400 1511.300 736.400 ;
      RECT 1513.260 1.400 1513.540 736.400 ;
      RECT 1515.500 1.400 1515.780 736.400 ;
      RECT 1517.740 1.400 1518.020 736.400 ;
      RECT 1519.980 1.400 1520.260 736.400 ;
      RECT 1522.220 1.400 1522.500 736.400 ;
      RECT 1524.460 1.400 1524.740 736.400 ;
      RECT 1526.700 1.400 1526.980 736.400 ;
      RECT 1528.940 1.400 1529.220 736.400 ;
      RECT 1531.180 1.400 1531.460 736.400 ;
      RECT 1533.420 1.400 1533.700 736.400 ;
      RECT 1535.660 1.400 1535.940 736.400 ;
      RECT 1537.900 1.400 1538.180 736.400 ;
      RECT 1540.140 1.400 1540.420 736.400 ;
      RECT 1542.380 1.400 1542.660 736.400 ;
      RECT 1544.620 1.400 1544.900 736.400 ;
      RECT 1546.860 1.400 1547.140 736.400 ;
      RECT 1549.100 1.400 1549.380 736.400 ;
      RECT 1551.340 1.400 1551.620 736.400 ;
      RECT 1553.580 1.400 1553.860 736.400 ;
      RECT 1555.820 1.400 1556.100 736.400 ;
      RECT 1558.060 1.400 1558.340 736.400 ;
      RECT 1560.300 1.400 1560.580 736.400 ;
      RECT 1562.540 1.400 1562.820 736.400 ;
      RECT 1564.780 1.400 1565.060 736.400 ;
      RECT 1567.020 1.400 1567.300 736.400 ;
      RECT 1569.260 1.400 1569.540 736.400 ;
      RECT 1571.500 1.400 1571.780 736.400 ;
      RECT 1573.740 1.400 1574.020 736.400 ;
      RECT 1575.980 1.400 1576.260 736.400 ;
      RECT 1578.220 1.400 1578.500 736.400 ;
      RECT 1580.460 1.400 1580.740 736.400 ;
      RECT 1582.700 1.400 1582.980 736.400 ;
      RECT 1584.940 1.400 1585.220 736.400 ;
      RECT 1587.180 1.400 1587.460 736.400 ;
      RECT 1589.420 1.400 1589.700 736.400 ;
      RECT 1591.660 1.400 1591.940 736.400 ;
      RECT 1593.900 1.400 1594.180 736.400 ;
      RECT 1596.140 1.400 1596.420 736.400 ;
      RECT 1598.380 1.400 1598.660 736.400 ;
      RECT 1600.620 1.400 1600.900 736.400 ;
      RECT 1602.860 1.400 1603.140 736.400 ;
      RECT 1605.100 1.400 1605.380 736.400 ;
      RECT 1607.340 1.400 1607.620 736.400 ;
      RECT 1609.580 1.400 1609.860 736.400 ;
      RECT 1611.820 1.400 1612.100 736.400 ;
      RECT 1614.060 1.400 1614.340 736.400 ;
      RECT 1616.300 1.400 1616.580 736.400 ;
      RECT 1618.540 1.400 1618.820 736.400 ;
      RECT 1620.780 1.400 1621.060 736.400 ;
      RECT 1623.020 1.400 1623.300 736.400 ;
      RECT 1625.260 1.400 1625.540 736.400 ;
      RECT 1627.500 1.400 1627.780 736.400 ;
      RECT 1629.740 1.400 1630.020 736.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 736.400 ;
      RECT 4.620 1.400 4.900 736.400 ;
      RECT 6.860 1.400 7.140 736.400 ;
      RECT 9.100 1.400 9.380 736.400 ;
      RECT 11.340 1.400 11.620 736.400 ;
      RECT 13.580 1.400 13.860 736.400 ;
      RECT 15.820 1.400 16.100 736.400 ;
      RECT 18.060 1.400 18.340 736.400 ;
      RECT 20.300 1.400 20.580 736.400 ;
      RECT 22.540 1.400 22.820 736.400 ;
      RECT 24.780 1.400 25.060 736.400 ;
      RECT 27.020 1.400 27.300 736.400 ;
      RECT 29.260 1.400 29.540 736.400 ;
      RECT 31.500 1.400 31.780 736.400 ;
      RECT 33.740 1.400 34.020 736.400 ;
      RECT 35.980 1.400 36.260 736.400 ;
      RECT 38.220 1.400 38.500 736.400 ;
      RECT 40.460 1.400 40.740 736.400 ;
      RECT 42.700 1.400 42.980 736.400 ;
      RECT 44.940 1.400 45.220 736.400 ;
      RECT 47.180 1.400 47.460 736.400 ;
      RECT 49.420 1.400 49.700 736.400 ;
      RECT 51.660 1.400 51.940 736.400 ;
      RECT 53.900 1.400 54.180 736.400 ;
      RECT 56.140 1.400 56.420 736.400 ;
      RECT 58.380 1.400 58.660 736.400 ;
      RECT 60.620 1.400 60.900 736.400 ;
      RECT 62.860 1.400 63.140 736.400 ;
      RECT 65.100 1.400 65.380 736.400 ;
      RECT 67.340 1.400 67.620 736.400 ;
      RECT 69.580 1.400 69.860 736.400 ;
      RECT 71.820 1.400 72.100 736.400 ;
      RECT 74.060 1.400 74.340 736.400 ;
      RECT 76.300 1.400 76.580 736.400 ;
      RECT 78.540 1.400 78.820 736.400 ;
      RECT 80.780 1.400 81.060 736.400 ;
      RECT 83.020 1.400 83.300 736.400 ;
      RECT 85.260 1.400 85.540 736.400 ;
      RECT 87.500 1.400 87.780 736.400 ;
      RECT 89.740 1.400 90.020 736.400 ;
      RECT 91.980 1.400 92.260 736.400 ;
      RECT 94.220 1.400 94.500 736.400 ;
      RECT 96.460 1.400 96.740 736.400 ;
      RECT 98.700 1.400 98.980 736.400 ;
      RECT 100.940 1.400 101.220 736.400 ;
      RECT 103.180 1.400 103.460 736.400 ;
      RECT 105.420 1.400 105.700 736.400 ;
      RECT 107.660 1.400 107.940 736.400 ;
      RECT 109.900 1.400 110.180 736.400 ;
      RECT 112.140 1.400 112.420 736.400 ;
      RECT 114.380 1.400 114.660 736.400 ;
      RECT 116.620 1.400 116.900 736.400 ;
      RECT 118.860 1.400 119.140 736.400 ;
      RECT 121.100 1.400 121.380 736.400 ;
      RECT 123.340 1.400 123.620 736.400 ;
      RECT 125.580 1.400 125.860 736.400 ;
      RECT 127.820 1.400 128.100 736.400 ;
      RECT 130.060 1.400 130.340 736.400 ;
      RECT 132.300 1.400 132.580 736.400 ;
      RECT 134.540 1.400 134.820 736.400 ;
      RECT 136.780 1.400 137.060 736.400 ;
      RECT 139.020 1.400 139.300 736.400 ;
      RECT 141.260 1.400 141.540 736.400 ;
      RECT 143.500 1.400 143.780 736.400 ;
      RECT 145.740 1.400 146.020 736.400 ;
      RECT 147.980 1.400 148.260 736.400 ;
      RECT 150.220 1.400 150.500 736.400 ;
      RECT 152.460 1.400 152.740 736.400 ;
      RECT 154.700 1.400 154.980 736.400 ;
      RECT 156.940 1.400 157.220 736.400 ;
      RECT 159.180 1.400 159.460 736.400 ;
      RECT 161.420 1.400 161.700 736.400 ;
      RECT 163.660 1.400 163.940 736.400 ;
      RECT 165.900 1.400 166.180 736.400 ;
      RECT 168.140 1.400 168.420 736.400 ;
      RECT 170.380 1.400 170.660 736.400 ;
      RECT 172.620 1.400 172.900 736.400 ;
      RECT 174.860 1.400 175.140 736.400 ;
      RECT 177.100 1.400 177.380 736.400 ;
      RECT 179.340 1.400 179.620 736.400 ;
      RECT 181.580 1.400 181.860 736.400 ;
      RECT 183.820 1.400 184.100 736.400 ;
      RECT 186.060 1.400 186.340 736.400 ;
      RECT 188.300 1.400 188.580 736.400 ;
      RECT 190.540 1.400 190.820 736.400 ;
      RECT 192.780 1.400 193.060 736.400 ;
      RECT 195.020 1.400 195.300 736.400 ;
      RECT 197.260 1.400 197.540 736.400 ;
      RECT 199.500 1.400 199.780 736.400 ;
      RECT 201.740 1.400 202.020 736.400 ;
      RECT 203.980 1.400 204.260 736.400 ;
      RECT 206.220 1.400 206.500 736.400 ;
      RECT 208.460 1.400 208.740 736.400 ;
      RECT 210.700 1.400 210.980 736.400 ;
      RECT 212.940 1.400 213.220 736.400 ;
      RECT 215.180 1.400 215.460 736.400 ;
      RECT 217.420 1.400 217.700 736.400 ;
      RECT 219.660 1.400 219.940 736.400 ;
      RECT 221.900 1.400 222.180 736.400 ;
      RECT 224.140 1.400 224.420 736.400 ;
      RECT 226.380 1.400 226.660 736.400 ;
      RECT 228.620 1.400 228.900 736.400 ;
      RECT 230.860 1.400 231.140 736.400 ;
      RECT 233.100 1.400 233.380 736.400 ;
      RECT 235.340 1.400 235.620 736.400 ;
      RECT 237.580 1.400 237.860 736.400 ;
      RECT 239.820 1.400 240.100 736.400 ;
      RECT 242.060 1.400 242.340 736.400 ;
      RECT 244.300 1.400 244.580 736.400 ;
      RECT 246.540 1.400 246.820 736.400 ;
      RECT 248.780 1.400 249.060 736.400 ;
      RECT 251.020 1.400 251.300 736.400 ;
      RECT 253.260 1.400 253.540 736.400 ;
      RECT 255.500 1.400 255.780 736.400 ;
      RECT 257.740 1.400 258.020 736.400 ;
      RECT 259.980 1.400 260.260 736.400 ;
      RECT 262.220 1.400 262.500 736.400 ;
      RECT 264.460 1.400 264.740 736.400 ;
      RECT 266.700 1.400 266.980 736.400 ;
      RECT 268.940 1.400 269.220 736.400 ;
      RECT 271.180 1.400 271.460 736.400 ;
      RECT 273.420 1.400 273.700 736.400 ;
      RECT 275.660 1.400 275.940 736.400 ;
      RECT 277.900 1.400 278.180 736.400 ;
      RECT 280.140 1.400 280.420 736.400 ;
      RECT 282.380 1.400 282.660 736.400 ;
      RECT 284.620 1.400 284.900 736.400 ;
      RECT 286.860 1.400 287.140 736.400 ;
      RECT 289.100 1.400 289.380 736.400 ;
      RECT 291.340 1.400 291.620 736.400 ;
      RECT 293.580 1.400 293.860 736.400 ;
      RECT 295.820 1.400 296.100 736.400 ;
      RECT 298.060 1.400 298.340 736.400 ;
      RECT 300.300 1.400 300.580 736.400 ;
      RECT 302.540 1.400 302.820 736.400 ;
      RECT 304.780 1.400 305.060 736.400 ;
      RECT 307.020 1.400 307.300 736.400 ;
      RECT 309.260 1.400 309.540 736.400 ;
      RECT 311.500 1.400 311.780 736.400 ;
      RECT 313.740 1.400 314.020 736.400 ;
      RECT 315.980 1.400 316.260 736.400 ;
      RECT 318.220 1.400 318.500 736.400 ;
      RECT 320.460 1.400 320.740 736.400 ;
      RECT 322.700 1.400 322.980 736.400 ;
      RECT 324.940 1.400 325.220 736.400 ;
      RECT 327.180 1.400 327.460 736.400 ;
      RECT 329.420 1.400 329.700 736.400 ;
      RECT 331.660 1.400 331.940 736.400 ;
      RECT 333.900 1.400 334.180 736.400 ;
      RECT 336.140 1.400 336.420 736.400 ;
      RECT 338.380 1.400 338.660 736.400 ;
      RECT 340.620 1.400 340.900 736.400 ;
      RECT 342.860 1.400 343.140 736.400 ;
      RECT 345.100 1.400 345.380 736.400 ;
      RECT 347.340 1.400 347.620 736.400 ;
      RECT 349.580 1.400 349.860 736.400 ;
      RECT 351.820 1.400 352.100 736.400 ;
      RECT 354.060 1.400 354.340 736.400 ;
      RECT 356.300 1.400 356.580 736.400 ;
      RECT 358.540 1.400 358.820 736.400 ;
      RECT 360.780 1.400 361.060 736.400 ;
      RECT 363.020 1.400 363.300 736.400 ;
      RECT 365.260 1.400 365.540 736.400 ;
      RECT 367.500 1.400 367.780 736.400 ;
      RECT 369.740 1.400 370.020 736.400 ;
      RECT 371.980 1.400 372.260 736.400 ;
      RECT 374.220 1.400 374.500 736.400 ;
      RECT 376.460 1.400 376.740 736.400 ;
      RECT 378.700 1.400 378.980 736.400 ;
      RECT 380.940 1.400 381.220 736.400 ;
      RECT 383.180 1.400 383.460 736.400 ;
      RECT 385.420 1.400 385.700 736.400 ;
      RECT 387.660 1.400 387.940 736.400 ;
      RECT 389.900 1.400 390.180 736.400 ;
      RECT 392.140 1.400 392.420 736.400 ;
      RECT 394.380 1.400 394.660 736.400 ;
      RECT 396.620 1.400 396.900 736.400 ;
      RECT 398.860 1.400 399.140 736.400 ;
      RECT 401.100 1.400 401.380 736.400 ;
      RECT 403.340 1.400 403.620 736.400 ;
      RECT 405.580 1.400 405.860 736.400 ;
      RECT 407.820 1.400 408.100 736.400 ;
      RECT 410.060 1.400 410.340 736.400 ;
      RECT 412.300 1.400 412.580 736.400 ;
      RECT 414.540 1.400 414.820 736.400 ;
      RECT 416.780 1.400 417.060 736.400 ;
      RECT 419.020 1.400 419.300 736.400 ;
      RECT 421.260 1.400 421.540 736.400 ;
      RECT 423.500 1.400 423.780 736.400 ;
      RECT 425.740 1.400 426.020 736.400 ;
      RECT 427.980 1.400 428.260 736.400 ;
      RECT 430.220 1.400 430.500 736.400 ;
      RECT 432.460 1.400 432.740 736.400 ;
      RECT 434.700 1.400 434.980 736.400 ;
      RECT 436.940 1.400 437.220 736.400 ;
      RECT 439.180 1.400 439.460 736.400 ;
      RECT 441.420 1.400 441.700 736.400 ;
      RECT 443.660 1.400 443.940 736.400 ;
      RECT 445.900 1.400 446.180 736.400 ;
      RECT 448.140 1.400 448.420 736.400 ;
      RECT 450.380 1.400 450.660 736.400 ;
      RECT 452.620 1.400 452.900 736.400 ;
      RECT 454.860 1.400 455.140 736.400 ;
      RECT 457.100 1.400 457.380 736.400 ;
      RECT 459.340 1.400 459.620 736.400 ;
      RECT 461.580 1.400 461.860 736.400 ;
      RECT 463.820 1.400 464.100 736.400 ;
      RECT 466.060 1.400 466.340 736.400 ;
      RECT 468.300 1.400 468.580 736.400 ;
      RECT 470.540 1.400 470.820 736.400 ;
      RECT 472.780 1.400 473.060 736.400 ;
      RECT 475.020 1.400 475.300 736.400 ;
      RECT 477.260 1.400 477.540 736.400 ;
      RECT 479.500 1.400 479.780 736.400 ;
      RECT 481.740 1.400 482.020 736.400 ;
      RECT 483.980 1.400 484.260 736.400 ;
      RECT 486.220 1.400 486.500 736.400 ;
      RECT 488.460 1.400 488.740 736.400 ;
      RECT 490.700 1.400 490.980 736.400 ;
      RECT 492.940 1.400 493.220 736.400 ;
      RECT 495.180 1.400 495.460 736.400 ;
      RECT 497.420 1.400 497.700 736.400 ;
      RECT 499.660 1.400 499.940 736.400 ;
      RECT 501.900 1.400 502.180 736.400 ;
      RECT 504.140 1.400 504.420 736.400 ;
      RECT 506.380 1.400 506.660 736.400 ;
      RECT 508.620 1.400 508.900 736.400 ;
      RECT 510.860 1.400 511.140 736.400 ;
      RECT 513.100 1.400 513.380 736.400 ;
      RECT 515.340 1.400 515.620 736.400 ;
      RECT 517.580 1.400 517.860 736.400 ;
      RECT 519.820 1.400 520.100 736.400 ;
      RECT 522.060 1.400 522.340 736.400 ;
      RECT 524.300 1.400 524.580 736.400 ;
      RECT 526.540 1.400 526.820 736.400 ;
      RECT 528.780 1.400 529.060 736.400 ;
      RECT 531.020 1.400 531.300 736.400 ;
      RECT 533.260 1.400 533.540 736.400 ;
      RECT 535.500 1.400 535.780 736.400 ;
      RECT 537.740 1.400 538.020 736.400 ;
      RECT 539.980 1.400 540.260 736.400 ;
      RECT 542.220 1.400 542.500 736.400 ;
      RECT 544.460 1.400 544.740 736.400 ;
      RECT 546.700 1.400 546.980 736.400 ;
      RECT 548.940 1.400 549.220 736.400 ;
      RECT 551.180 1.400 551.460 736.400 ;
      RECT 553.420 1.400 553.700 736.400 ;
      RECT 555.660 1.400 555.940 736.400 ;
      RECT 557.900 1.400 558.180 736.400 ;
      RECT 560.140 1.400 560.420 736.400 ;
      RECT 562.380 1.400 562.660 736.400 ;
      RECT 564.620 1.400 564.900 736.400 ;
      RECT 566.860 1.400 567.140 736.400 ;
      RECT 569.100 1.400 569.380 736.400 ;
      RECT 571.340 1.400 571.620 736.400 ;
      RECT 573.580 1.400 573.860 736.400 ;
      RECT 575.820 1.400 576.100 736.400 ;
      RECT 578.060 1.400 578.340 736.400 ;
      RECT 580.300 1.400 580.580 736.400 ;
      RECT 582.540 1.400 582.820 736.400 ;
      RECT 584.780 1.400 585.060 736.400 ;
      RECT 587.020 1.400 587.300 736.400 ;
      RECT 589.260 1.400 589.540 736.400 ;
      RECT 591.500 1.400 591.780 736.400 ;
      RECT 593.740 1.400 594.020 736.400 ;
      RECT 595.980 1.400 596.260 736.400 ;
      RECT 598.220 1.400 598.500 736.400 ;
      RECT 600.460 1.400 600.740 736.400 ;
      RECT 602.700 1.400 602.980 736.400 ;
      RECT 604.940 1.400 605.220 736.400 ;
      RECT 607.180 1.400 607.460 736.400 ;
      RECT 609.420 1.400 609.700 736.400 ;
      RECT 611.660 1.400 611.940 736.400 ;
      RECT 613.900 1.400 614.180 736.400 ;
      RECT 616.140 1.400 616.420 736.400 ;
      RECT 618.380 1.400 618.660 736.400 ;
      RECT 620.620 1.400 620.900 736.400 ;
      RECT 622.860 1.400 623.140 736.400 ;
      RECT 625.100 1.400 625.380 736.400 ;
      RECT 627.340 1.400 627.620 736.400 ;
      RECT 629.580 1.400 629.860 736.400 ;
      RECT 631.820 1.400 632.100 736.400 ;
      RECT 634.060 1.400 634.340 736.400 ;
      RECT 636.300 1.400 636.580 736.400 ;
      RECT 638.540 1.400 638.820 736.400 ;
      RECT 640.780 1.400 641.060 736.400 ;
      RECT 643.020 1.400 643.300 736.400 ;
      RECT 645.260 1.400 645.540 736.400 ;
      RECT 647.500 1.400 647.780 736.400 ;
      RECT 649.740 1.400 650.020 736.400 ;
      RECT 651.980 1.400 652.260 736.400 ;
      RECT 654.220 1.400 654.500 736.400 ;
      RECT 656.460 1.400 656.740 736.400 ;
      RECT 658.700 1.400 658.980 736.400 ;
      RECT 660.940 1.400 661.220 736.400 ;
      RECT 663.180 1.400 663.460 736.400 ;
      RECT 665.420 1.400 665.700 736.400 ;
      RECT 667.660 1.400 667.940 736.400 ;
      RECT 669.900 1.400 670.180 736.400 ;
      RECT 672.140 1.400 672.420 736.400 ;
      RECT 674.380 1.400 674.660 736.400 ;
      RECT 676.620 1.400 676.900 736.400 ;
      RECT 678.860 1.400 679.140 736.400 ;
      RECT 681.100 1.400 681.380 736.400 ;
      RECT 683.340 1.400 683.620 736.400 ;
      RECT 685.580 1.400 685.860 736.400 ;
      RECT 687.820 1.400 688.100 736.400 ;
      RECT 690.060 1.400 690.340 736.400 ;
      RECT 692.300 1.400 692.580 736.400 ;
      RECT 694.540 1.400 694.820 736.400 ;
      RECT 696.780 1.400 697.060 736.400 ;
      RECT 699.020 1.400 699.300 736.400 ;
      RECT 701.260 1.400 701.540 736.400 ;
      RECT 703.500 1.400 703.780 736.400 ;
      RECT 705.740 1.400 706.020 736.400 ;
      RECT 707.980 1.400 708.260 736.400 ;
      RECT 710.220 1.400 710.500 736.400 ;
      RECT 712.460 1.400 712.740 736.400 ;
      RECT 714.700 1.400 714.980 736.400 ;
      RECT 716.940 1.400 717.220 736.400 ;
      RECT 719.180 1.400 719.460 736.400 ;
      RECT 721.420 1.400 721.700 736.400 ;
      RECT 723.660 1.400 723.940 736.400 ;
      RECT 725.900 1.400 726.180 736.400 ;
      RECT 728.140 1.400 728.420 736.400 ;
      RECT 730.380 1.400 730.660 736.400 ;
      RECT 732.620 1.400 732.900 736.400 ;
      RECT 734.860 1.400 735.140 736.400 ;
      RECT 737.100 1.400 737.380 736.400 ;
      RECT 739.340 1.400 739.620 736.400 ;
      RECT 741.580 1.400 741.860 736.400 ;
      RECT 743.820 1.400 744.100 736.400 ;
      RECT 746.060 1.400 746.340 736.400 ;
      RECT 748.300 1.400 748.580 736.400 ;
      RECT 750.540 1.400 750.820 736.400 ;
      RECT 752.780 1.400 753.060 736.400 ;
      RECT 755.020 1.400 755.300 736.400 ;
      RECT 757.260 1.400 757.540 736.400 ;
      RECT 759.500 1.400 759.780 736.400 ;
      RECT 761.740 1.400 762.020 736.400 ;
      RECT 763.980 1.400 764.260 736.400 ;
      RECT 766.220 1.400 766.500 736.400 ;
      RECT 768.460 1.400 768.740 736.400 ;
      RECT 770.700 1.400 770.980 736.400 ;
      RECT 772.940 1.400 773.220 736.400 ;
      RECT 775.180 1.400 775.460 736.400 ;
      RECT 777.420 1.400 777.700 736.400 ;
      RECT 779.660 1.400 779.940 736.400 ;
      RECT 781.900 1.400 782.180 736.400 ;
      RECT 784.140 1.400 784.420 736.400 ;
      RECT 786.380 1.400 786.660 736.400 ;
      RECT 788.620 1.400 788.900 736.400 ;
      RECT 790.860 1.400 791.140 736.400 ;
      RECT 793.100 1.400 793.380 736.400 ;
      RECT 795.340 1.400 795.620 736.400 ;
      RECT 797.580 1.400 797.860 736.400 ;
      RECT 799.820 1.400 800.100 736.400 ;
      RECT 802.060 1.400 802.340 736.400 ;
      RECT 804.300 1.400 804.580 736.400 ;
      RECT 806.540 1.400 806.820 736.400 ;
      RECT 808.780 1.400 809.060 736.400 ;
      RECT 811.020 1.400 811.300 736.400 ;
      RECT 813.260 1.400 813.540 736.400 ;
      RECT 815.500 1.400 815.780 736.400 ;
      RECT 817.740 1.400 818.020 736.400 ;
      RECT 819.980 1.400 820.260 736.400 ;
      RECT 822.220 1.400 822.500 736.400 ;
      RECT 824.460 1.400 824.740 736.400 ;
      RECT 826.700 1.400 826.980 736.400 ;
      RECT 828.940 1.400 829.220 736.400 ;
      RECT 831.180 1.400 831.460 736.400 ;
      RECT 833.420 1.400 833.700 736.400 ;
      RECT 835.660 1.400 835.940 736.400 ;
      RECT 837.900 1.400 838.180 736.400 ;
      RECT 840.140 1.400 840.420 736.400 ;
      RECT 842.380 1.400 842.660 736.400 ;
      RECT 844.620 1.400 844.900 736.400 ;
      RECT 846.860 1.400 847.140 736.400 ;
      RECT 849.100 1.400 849.380 736.400 ;
      RECT 851.340 1.400 851.620 736.400 ;
      RECT 853.580 1.400 853.860 736.400 ;
      RECT 855.820 1.400 856.100 736.400 ;
      RECT 858.060 1.400 858.340 736.400 ;
      RECT 860.300 1.400 860.580 736.400 ;
      RECT 862.540 1.400 862.820 736.400 ;
      RECT 864.780 1.400 865.060 736.400 ;
      RECT 867.020 1.400 867.300 736.400 ;
      RECT 869.260 1.400 869.540 736.400 ;
      RECT 871.500 1.400 871.780 736.400 ;
      RECT 873.740 1.400 874.020 736.400 ;
      RECT 875.980 1.400 876.260 736.400 ;
      RECT 878.220 1.400 878.500 736.400 ;
      RECT 880.460 1.400 880.740 736.400 ;
      RECT 882.700 1.400 882.980 736.400 ;
      RECT 884.940 1.400 885.220 736.400 ;
      RECT 887.180 1.400 887.460 736.400 ;
      RECT 889.420 1.400 889.700 736.400 ;
      RECT 891.660 1.400 891.940 736.400 ;
      RECT 893.900 1.400 894.180 736.400 ;
      RECT 896.140 1.400 896.420 736.400 ;
      RECT 898.380 1.400 898.660 736.400 ;
      RECT 900.620 1.400 900.900 736.400 ;
      RECT 902.860 1.400 903.140 736.400 ;
      RECT 905.100 1.400 905.380 736.400 ;
      RECT 907.340 1.400 907.620 736.400 ;
      RECT 909.580 1.400 909.860 736.400 ;
      RECT 911.820 1.400 912.100 736.400 ;
      RECT 914.060 1.400 914.340 736.400 ;
      RECT 916.300 1.400 916.580 736.400 ;
      RECT 918.540 1.400 918.820 736.400 ;
      RECT 920.780 1.400 921.060 736.400 ;
      RECT 923.020 1.400 923.300 736.400 ;
      RECT 925.260 1.400 925.540 736.400 ;
      RECT 927.500 1.400 927.780 736.400 ;
      RECT 929.740 1.400 930.020 736.400 ;
      RECT 931.980 1.400 932.260 736.400 ;
      RECT 934.220 1.400 934.500 736.400 ;
      RECT 936.460 1.400 936.740 736.400 ;
      RECT 938.700 1.400 938.980 736.400 ;
      RECT 940.940 1.400 941.220 736.400 ;
      RECT 943.180 1.400 943.460 736.400 ;
      RECT 945.420 1.400 945.700 736.400 ;
      RECT 947.660 1.400 947.940 736.400 ;
      RECT 949.900 1.400 950.180 736.400 ;
      RECT 952.140 1.400 952.420 736.400 ;
      RECT 954.380 1.400 954.660 736.400 ;
      RECT 956.620 1.400 956.900 736.400 ;
      RECT 958.860 1.400 959.140 736.400 ;
      RECT 961.100 1.400 961.380 736.400 ;
      RECT 963.340 1.400 963.620 736.400 ;
      RECT 965.580 1.400 965.860 736.400 ;
      RECT 967.820 1.400 968.100 736.400 ;
      RECT 970.060 1.400 970.340 736.400 ;
      RECT 972.300 1.400 972.580 736.400 ;
      RECT 974.540 1.400 974.820 736.400 ;
      RECT 976.780 1.400 977.060 736.400 ;
      RECT 979.020 1.400 979.300 736.400 ;
      RECT 981.260 1.400 981.540 736.400 ;
      RECT 983.500 1.400 983.780 736.400 ;
      RECT 985.740 1.400 986.020 736.400 ;
      RECT 987.980 1.400 988.260 736.400 ;
      RECT 990.220 1.400 990.500 736.400 ;
      RECT 992.460 1.400 992.740 736.400 ;
      RECT 994.700 1.400 994.980 736.400 ;
      RECT 996.940 1.400 997.220 736.400 ;
      RECT 999.180 1.400 999.460 736.400 ;
      RECT 1001.420 1.400 1001.700 736.400 ;
      RECT 1003.660 1.400 1003.940 736.400 ;
      RECT 1005.900 1.400 1006.180 736.400 ;
      RECT 1008.140 1.400 1008.420 736.400 ;
      RECT 1010.380 1.400 1010.660 736.400 ;
      RECT 1012.620 1.400 1012.900 736.400 ;
      RECT 1014.860 1.400 1015.140 736.400 ;
      RECT 1017.100 1.400 1017.380 736.400 ;
      RECT 1019.340 1.400 1019.620 736.400 ;
      RECT 1021.580 1.400 1021.860 736.400 ;
      RECT 1023.820 1.400 1024.100 736.400 ;
      RECT 1026.060 1.400 1026.340 736.400 ;
      RECT 1028.300 1.400 1028.580 736.400 ;
      RECT 1030.540 1.400 1030.820 736.400 ;
      RECT 1032.780 1.400 1033.060 736.400 ;
      RECT 1035.020 1.400 1035.300 736.400 ;
      RECT 1037.260 1.400 1037.540 736.400 ;
      RECT 1039.500 1.400 1039.780 736.400 ;
      RECT 1041.740 1.400 1042.020 736.400 ;
      RECT 1043.980 1.400 1044.260 736.400 ;
      RECT 1046.220 1.400 1046.500 736.400 ;
      RECT 1048.460 1.400 1048.740 736.400 ;
      RECT 1050.700 1.400 1050.980 736.400 ;
      RECT 1052.940 1.400 1053.220 736.400 ;
      RECT 1055.180 1.400 1055.460 736.400 ;
      RECT 1057.420 1.400 1057.700 736.400 ;
      RECT 1059.660 1.400 1059.940 736.400 ;
      RECT 1061.900 1.400 1062.180 736.400 ;
      RECT 1064.140 1.400 1064.420 736.400 ;
      RECT 1066.380 1.400 1066.660 736.400 ;
      RECT 1068.620 1.400 1068.900 736.400 ;
      RECT 1070.860 1.400 1071.140 736.400 ;
      RECT 1073.100 1.400 1073.380 736.400 ;
      RECT 1075.340 1.400 1075.620 736.400 ;
      RECT 1077.580 1.400 1077.860 736.400 ;
      RECT 1079.820 1.400 1080.100 736.400 ;
      RECT 1082.060 1.400 1082.340 736.400 ;
      RECT 1084.300 1.400 1084.580 736.400 ;
      RECT 1086.540 1.400 1086.820 736.400 ;
      RECT 1088.780 1.400 1089.060 736.400 ;
      RECT 1091.020 1.400 1091.300 736.400 ;
      RECT 1093.260 1.400 1093.540 736.400 ;
      RECT 1095.500 1.400 1095.780 736.400 ;
      RECT 1097.740 1.400 1098.020 736.400 ;
      RECT 1099.980 1.400 1100.260 736.400 ;
      RECT 1102.220 1.400 1102.500 736.400 ;
      RECT 1104.460 1.400 1104.740 736.400 ;
      RECT 1106.700 1.400 1106.980 736.400 ;
      RECT 1108.940 1.400 1109.220 736.400 ;
      RECT 1111.180 1.400 1111.460 736.400 ;
      RECT 1113.420 1.400 1113.700 736.400 ;
      RECT 1115.660 1.400 1115.940 736.400 ;
      RECT 1117.900 1.400 1118.180 736.400 ;
      RECT 1120.140 1.400 1120.420 736.400 ;
      RECT 1122.380 1.400 1122.660 736.400 ;
      RECT 1124.620 1.400 1124.900 736.400 ;
      RECT 1126.860 1.400 1127.140 736.400 ;
      RECT 1129.100 1.400 1129.380 736.400 ;
      RECT 1131.340 1.400 1131.620 736.400 ;
      RECT 1133.580 1.400 1133.860 736.400 ;
      RECT 1135.820 1.400 1136.100 736.400 ;
      RECT 1138.060 1.400 1138.340 736.400 ;
      RECT 1140.300 1.400 1140.580 736.400 ;
      RECT 1142.540 1.400 1142.820 736.400 ;
      RECT 1144.780 1.400 1145.060 736.400 ;
      RECT 1147.020 1.400 1147.300 736.400 ;
      RECT 1149.260 1.400 1149.540 736.400 ;
      RECT 1151.500 1.400 1151.780 736.400 ;
      RECT 1153.740 1.400 1154.020 736.400 ;
      RECT 1155.980 1.400 1156.260 736.400 ;
      RECT 1158.220 1.400 1158.500 736.400 ;
      RECT 1160.460 1.400 1160.740 736.400 ;
      RECT 1162.700 1.400 1162.980 736.400 ;
      RECT 1164.940 1.400 1165.220 736.400 ;
      RECT 1167.180 1.400 1167.460 736.400 ;
      RECT 1169.420 1.400 1169.700 736.400 ;
      RECT 1171.660 1.400 1171.940 736.400 ;
      RECT 1173.900 1.400 1174.180 736.400 ;
      RECT 1176.140 1.400 1176.420 736.400 ;
      RECT 1178.380 1.400 1178.660 736.400 ;
      RECT 1180.620 1.400 1180.900 736.400 ;
      RECT 1182.860 1.400 1183.140 736.400 ;
      RECT 1185.100 1.400 1185.380 736.400 ;
      RECT 1187.340 1.400 1187.620 736.400 ;
      RECT 1189.580 1.400 1189.860 736.400 ;
      RECT 1191.820 1.400 1192.100 736.400 ;
      RECT 1194.060 1.400 1194.340 736.400 ;
      RECT 1196.300 1.400 1196.580 736.400 ;
      RECT 1198.540 1.400 1198.820 736.400 ;
      RECT 1200.780 1.400 1201.060 736.400 ;
      RECT 1203.020 1.400 1203.300 736.400 ;
      RECT 1205.260 1.400 1205.540 736.400 ;
      RECT 1207.500 1.400 1207.780 736.400 ;
      RECT 1209.740 1.400 1210.020 736.400 ;
      RECT 1211.980 1.400 1212.260 736.400 ;
      RECT 1214.220 1.400 1214.500 736.400 ;
      RECT 1216.460 1.400 1216.740 736.400 ;
      RECT 1218.700 1.400 1218.980 736.400 ;
      RECT 1220.940 1.400 1221.220 736.400 ;
      RECT 1223.180 1.400 1223.460 736.400 ;
      RECT 1225.420 1.400 1225.700 736.400 ;
      RECT 1227.660 1.400 1227.940 736.400 ;
      RECT 1229.900 1.400 1230.180 736.400 ;
      RECT 1232.140 1.400 1232.420 736.400 ;
      RECT 1234.380 1.400 1234.660 736.400 ;
      RECT 1236.620 1.400 1236.900 736.400 ;
      RECT 1238.860 1.400 1239.140 736.400 ;
      RECT 1241.100 1.400 1241.380 736.400 ;
      RECT 1243.340 1.400 1243.620 736.400 ;
      RECT 1245.580 1.400 1245.860 736.400 ;
      RECT 1247.820 1.400 1248.100 736.400 ;
      RECT 1250.060 1.400 1250.340 736.400 ;
      RECT 1252.300 1.400 1252.580 736.400 ;
      RECT 1254.540 1.400 1254.820 736.400 ;
      RECT 1256.780 1.400 1257.060 736.400 ;
      RECT 1259.020 1.400 1259.300 736.400 ;
      RECT 1261.260 1.400 1261.540 736.400 ;
      RECT 1263.500 1.400 1263.780 736.400 ;
      RECT 1265.740 1.400 1266.020 736.400 ;
      RECT 1267.980 1.400 1268.260 736.400 ;
      RECT 1270.220 1.400 1270.500 736.400 ;
      RECT 1272.460 1.400 1272.740 736.400 ;
      RECT 1274.700 1.400 1274.980 736.400 ;
      RECT 1276.940 1.400 1277.220 736.400 ;
      RECT 1279.180 1.400 1279.460 736.400 ;
      RECT 1281.420 1.400 1281.700 736.400 ;
      RECT 1283.660 1.400 1283.940 736.400 ;
      RECT 1285.900 1.400 1286.180 736.400 ;
      RECT 1288.140 1.400 1288.420 736.400 ;
      RECT 1290.380 1.400 1290.660 736.400 ;
      RECT 1292.620 1.400 1292.900 736.400 ;
      RECT 1294.860 1.400 1295.140 736.400 ;
      RECT 1297.100 1.400 1297.380 736.400 ;
      RECT 1299.340 1.400 1299.620 736.400 ;
      RECT 1301.580 1.400 1301.860 736.400 ;
      RECT 1303.820 1.400 1304.100 736.400 ;
      RECT 1306.060 1.400 1306.340 736.400 ;
      RECT 1308.300 1.400 1308.580 736.400 ;
      RECT 1310.540 1.400 1310.820 736.400 ;
      RECT 1312.780 1.400 1313.060 736.400 ;
      RECT 1315.020 1.400 1315.300 736.400 ;
      RECT 1317.260 1.400 1317.540 736.400 ;
      RECT 1319.500 1.400 1319.780 736.400 ;
      RECT 1321.740 1.400 1322.020 736.400 ;
      RECT 1323.980 1.400 1324.260 736.400 ;
      RECT 1326.220 1.400 1326.500 736.400 ;
      RECT 1328.460 1.400 1328.740 736.400 ;
      RECT 1330.700 1.400 1330.980 736.400 ;
      RECT 1332.940 1.400 1333.220 736.400 ;
      RECT 1335.180 1.400 1335.460 736.400 ;
      RECT 1337.420 1.400 1337.700 736.400 ;
      RECT 1339.660 1.400 1339.940 736.400 ;
      RECT 1341.900 1.400 1342.180 736.400 ;
      RECT 1344.140 1.400 1344.420 736.400 ;
      RECT 1346.380 1.400 1346.660 736.400 ;
      RECT 1348.620 1.400 1348.900 736.400 ;
      RECT 1350.860 1.400 1351.140 736.400 ;
      RECT 1353.100 1.400 1353.380 736.400 ;
      RECT 1355.340 1.400 1355.620 736.400 ;
      RECT 1357.580 1.400 1357.860 736.400 ;
      RECT 1359.820 1.400 1360.100 736.400 ;
      RECT 1362.060 1.400 1362.340 736.400 ;
      RECT 1364.300 1.400 1364.580 736.400 ;
      RECT 1366.540 1.400 1366.820 736.400 ;
      RECT 1368.780 1.400 1369.060 736.400 ;
      RECT 1371.020 1.400 1371.300 736.400 ;
      RECT 1373.260 1.400 1373.540 736.400 ;
      RECT 1375.500 1.400 1375.780 736.400 ;
      RECT 1377.740 1.400 1378.020 736.400 ;
      RECT 1379.980 1.400 1380.260 736.400 ;
      RECT 1382.220 1.400 1382.500 736.400 ;
      RECT 1384.460 1.400 1384.740 736.400 ;
      RECT 1386.700 1.400 1386.980 736.400 ;
      RECT 1388.940 1.400 1389.220 736.400 ;
      RECT 1391.180 1.400 1391.460 736.400 ;
      RECT 1393.420 1.400 1393.700 736.400 ;
      RECT 1395.660 1.400 1395.940 736.400 ;
      RECT 1397.900 1.400 1398.180 736.400 ;
      RECT 1400.140 1.400 1400.420 736.400 ;
      RECT 1402.380 1.400 1402.660 736.400 ;
      RECT 1404.620 1.400 1404.900 736.400 ;
      RECT 1406.860 1.400 1407.140 736.400 ;
      RECT 1409.100 1.400 1409.380 736.400 ;
      RECT 1411.340 1.400 1411.620 736.400 ;
      RECT 1413.580 1.400 1413.860 736.400 ;
      RECT 1415.820 1.400 1416.100 736.400 ;
      RECT 1418.060 1.400 1418.340 736.400 ;
      RECT 1420.300 1.400 1420.580 736.400 ;
      RECT 1422.540 1.400 1422.820 736.400 ;
      RECT 1424.780 1.400 1425.060 736.400 ;
      RECT 1427.020 1.400 1427.300 736.400 ;
      RECT 1429.260 1.400 1429.540 736.400 ;
      RECT 1431.500 1.400 1431.780 736.400 ;
      RECT 1433.740 1.400 1434.020 736.400 ;
      RECT 1435.980 1.400 1436.260 736.400 ;
      RECT 1438.220 1.400 1438.500 736.400 ;
      RECT 1440.460 1.400 1440.740 736.400 ;
      RECT 1442.700 1.400 1442.980 736.400 ;
      RECT 1444.940 1.400 1445.220 736.400 ;
      RECT 1447.180 1.400 1447.460 736.400 ;
      RECT 1449.420 1.400 1449.700 736.400 ;
      RECT 1451.660 1.400 1451.940 736.400 ;
      RECT 1453.900 1.400 1454.180 736.400 ;
      RECT 1456.140 1.400 1456.420 736.400 ;
      RECT 1458.380 1.400 1458.660 736.400 ;
      RECT 1460.620 1.400 1460.900 736.400 ;
      RECT 1462.860 1.400 1463.140 736.400 ;
      RECT 1465.100 1.400 1465.380 736.400 ;
      RECT 1467.340 1.400 1467.620 736.400 ;
      RECT 1469.580 1.400 1469.860 736.400 ;
      RECT 1471.820 1.400 1472.100 736.400 ;
      RECT 1474.060 1.400 1474.340 736.400 ;
      RECT 1476.300 1.400 1476.580 736.400 ;
      RECT 1478.540 1.400 1478.820 736.400 ;
      RECT 1480.780 1.400 1481.060 736.400 ;
      RECT 1483.020 1.400 1483.300 736.400 ;
      RECT 1485.260 1.400 1485.540 736.400 ;
      RECT 1487.500 1.400 1487.780 736.400 ;
      RECT 1489.740 1.400 1490.020 736.400 ;
      RECT 1491.980 1.400 1492.260 736.400 ;
      RECT 1494.220 1.400 1494.500 736.400 ;
      RECT 1496.460 1.400 1496.740 736.400 ;
      RECT 1498.700 1.400 1498.980 736.400 ;
      RECT 1500.940 1.400 1501.220 736.400 ;
      RECT 1503.180 1.400 1503.460 736.400 ;
      RECT 1505.420 1.400 1505.700 736.400 ;
      RECT 1507.660 1.400 1507.940 736.400 ;
      RECT 1509.900 1.400 1510.180 736.400 ;
      RECT 1512.140 1.400 1512.420 736.400 ;
      RECT 1514.380 1.400 1514.660 736.400 ;
      RECT 1516.620 1.400 1516.900 736.400 ;
      RECT 1518.860 1.400 1519.140 736.400 ;
      RECT 1521.100 1.400 1521.380 736.400 ;
      RECT 1523.340 1.400 1523.620 736.400 ;
      RECT 1525.580 1.400 1525.860 736.400 ;
      RECT 1527.820 1.400 1528.100 736.400 ;
      RECT 1530.060 1.400 1530.340 736.400 ;
      RECT 1532.300 1.400 1532.580 736.400 ;
      RECT 1534.540 1.400 1534.820 736.400 ;
      RECT 1536.780 1.400 1537.060 736.400 ;
      RECT 1539.020 1.400 1539.300 736.400 ;
      RECT 1541.260 1.400 1541.540 736.400 ;
      RECT 1543.500 1.400 1543.780 736.400 ;
      RECT 1545.740 1.400 1546.020 736.400 ;
      RECT 1547.980 1.400 1548.260 736.400 ;
      RECT 1550.220 1.400 1550.500 736.400 ;
      RECT 1552.460 1.400 1552.740 736.400 ;
      RECT 1554.700 1.400 1554.980 736.400 ;
      RECT 1556.940 1.400 1557.220 736.400 ;
      RECT 1559.180 1.400 1559.460 736.400 ;
      RECT 1561.420 1.400 1561.700 736.400 ;
      RECT 1563.660 1.400 1563.940 736.400 ;
      RECT 1565.900 1.400 1566.180 736.400 ;
      RECT 1568.140 1.400 1568.420 736.400 ;
      RECT 1570.380 1.400 1570.660 736.400 ;
      RECT 1572.620 1.400 1572.900 736.400 ;
      RECT 1574.860 1.400 1575.140 736.400 ;
      RECT 1577.100 1.400 1577.380 736.400 ;
      RECT 1579.340 1.400 1579.620 736.400 ;
      RECT 1581.580 1.400 1581.860 736.400 ;
      RECT 1583.820 1.400 1584.100 736.400 ;
      RECT 1586.060 1.400 1586.340 736.400 ;
      RECT 1588.300 1.400 1588.580 736.400 ;
      RECT 1590.540 1.400 1590.820 736.400 ;
      RECT 1592.780 1.400 1593.060 736.400 ;
      RECT 1595.020 1.400 1595.300 736.400 ;
      RECT 1597.260 1.400 1597.540 736.400 ;
      RECT 1599.500 1.400 1599.780 736.400 ;
      RECT 1601.740 1.400 1602.020 736.400 ;
      RECT 1603.980 1.400 1604.260 736.400 ;
      RECT 1606.220 1.400 1606.500 736.400 ;
      RECT 1608.460 1.400 1608.740 736.400 ;
      RECT 1610.700 1.400 1610.980 736.400 ;
      RECT 1612.940 1.400 1613.220 736.400 ;
      RECT 1615.180 1.400 1615.460 736.400 ;
      RECT 1617.420 1.400 1617.700 736.400 ;
      RECT 1619.660 1.400 1619.940 736.400 ;
      RECT 1621.900 1.400 1622.180 736.400 ;
      RECT 1624.140 1.400 1624.420 736.400 ;
      RECT 1626.380 1.400 1626.660 736.400 ;
      RECT 1628.620 1.400 1628.900 736.400 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 1631.530 737.800 ;
    LAYER metal2 ;
    RECT 0 0 1631.530 737.800 ;
    LAYER metal3 ;
    RECT 0.070 0 1631.530 737.800 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.205 ;
    RECT 0 2.275 0.070 3.045 ;
    RECT 0 3.115 0.070 3.885 ;
    RECT 0 3.955 0.070 4.725 ;
    RECT 0 4.795 0.070 5.565 ;
    RECT 0 5.635 0.070 6.405 ;
    RECT 0 6.475 0.070 7.245 ;
    RECT 0 7.315 0.070 8.085 ;
    RECT 0 8.155 0.070 8.925 ;
    RECT 0 8.995 0.070 9.765 ;
    RECT 0 9.835 0.070 10.605 ;
    RECT 0 10.675 0.070 11.445 ;
    RECT 0 11.515 0.070 12.285 ;
    RECT 0 12.355 0.070 13.125 ;
    RECT 0 13.195 0.070 13.965 ;
    RECT 0 14.035 0.070 14.805 ;
    RECT 0 14.875 0.070 15.645 ;
    RECT 0 15.715 0.070 16.485 ;
    RECT 0 16.555 0.070 17.325 ;
    RECT 0 17.395 0.070 18.165 ;
    RECT 0 18.235 0.070 19.005 ;
    RECT 0 19.075 0.070 19.845 ;
    RECT 0 19.915 0.070 20.685 ;
    RECT 0 20.755 0.070 21.525 ;
    RECT 0 21.595 0.070 22.365 ;
    RECT 0 22.435 0.070 23.205 ;
    RECT 0 23.275 0.070 24.045 ;
    RECT 0 24.115 0.070 24.885 ;
    RECT 0 24.955 0.070 25.725 ;
    RECT 0 25.795 0.070 26.565 ;
    RECT 0 26.635 0.070 27.405 ;
    RECT 0 27.475 0.070 28.245 ;
    RECT 0 28.315 0.070 29.085 ;
    RECT 0 29.155 0.070 29.925 ;
    RECT 0 29.995 0.070 30.765 ;
    RECT 0 30.835 0.070 31.605 ;
    RECT 0 31.675 0.070 32.445 ;
    RECT 0 32.515 0.070 33.285 ;
    RECT 0 33.355 0.070 34.125 ;
    RECT 0 34.195 0.070 34.965 ;
    RECT 0 35.035 0.070 35.805 ;
    RECT 0 35.875 0.070 36.645 ;
    RECT 0 36.715 0.070 37.485 ;
    RECT 0 37.555 0.070 38.325 ;
    RECT 0 38.395 0.070 39.165 ;
    RECT 0 39.235 0.070 40.005 ;
    RECT 0 40.075 0.070 40.845 ;
    RECT 0 40.915 0.070 41.685 ;
    RECT 0 41.755 0.070 42.525 ;
    RECT 0 42.595 0.070 43.365 ;
    RECT 0 43.435 0.070 44.205 ;
    RECT 0 44.275 0.070 45.045 ;
    RECT 0 45.115 0.070 45.885 ;
    RECT 0 45.955 0.070 46.725 ;
    RECT 0 46.795 0.070 47.565 ;
    RECT 0 47.635 0.070 48.405 ;
    RECT 0 48.475 0.070 49.245 ;
    RECT 0 49.315 0.070 50.085 ;
    RECT 0 50.155 0.070 50.925 ;
    RECT 0 50.995 0.070 51.765 ;
    RECT 0 51.835 0.070 52.605 ;
    RECT 0 52.675 0.070 53.445 ;
    RECT 0 53.515 0.070 54.285 ;
    RECT 0 54.355 0.070 55.125 ;
    RECT 0 55.195 0.070 55.965 ;
    RECT 0 56.035 0.070 56.805 ;
    RECT 0 56.875 0.070 57.645 ;
    RECT 0 57.715 0.070 58.485 ;
    RECT 0 58.555 0.070 59.325 ;
    RECT 0 59.395 0.070 60.165 ;
    RECT 0 60.235 0.070 61.005 ;
    RECT 0 61.075 0.070 61.845 ;
    RECT 0 61.915 0.070 62.685 ;
    RECT 0 62.755 0.070 63.525 ;
    RECT 0 63.595 0.070 64.365 ;
    RECT 0 64.435 0.070 65.205 ;
    RECT 0 65.275 0.070 66.045 ;
    RECT 0 66.115 0.070 66.885 ;
    RECT 0 66.955 0.070 67.725 ;
    RECT 0 67.795 0.070 68.565 ;
    RECT 0 68.635 0.070 69.405 ;
    RECT 0 69.475 0.070 70.245 ;
    RECT 0 70.315 0.070 71.085 ;
    RECT 0 71.155 0.070 71.925 ;
    RECT 0 71.995 0.070 72.765 ;
    RECT 0 72.835 0.070 73.605 ;
    RECT 0 73.675 0.070 74.445 ;
    RECT 0 74.515 0.070 75.285 ;
    RECT 0 75.355 0.070 76.125 ;
    RECT 0 76.195 0.070 76.965 ;
    RECT 0 77.035 0.070 77.805 ;
    RECT 0 77.875 0.070 78.645 ;
    RECT 0 78.715 0.070 79.485 ;
    RECT 0 79.555 0.070 80.325 ;
    RECT 0 80.395 0.070 81.165 ;
    RECT 0 81.235 0.070 82.005 ;
    RECT 0 82.075 0.070 82.845 ;
    RECT 0 82.915 0.070 83.685 ;
    RECT 0 83.755 0.070 84.525 ;
    RECT 0 84.595 0.070 85.365 ;
    RECT 0 85.435 0.070 86.205 ;
    RECT 0 86.275 0.070 87.045 ;
    RECT 0 87.115 0.070 87.885 ;
    RECT 0 87.955 0.070 88.725 ;
    RECT 0 88.795 0.070 89.565 ;
    RECT 0 89.635 0.070 90.405 ;
    RECT 0 90.475 0.070 91.245 ;
    RECT 0 91.315 0.070 92.085 ;
    RECT 0 92.155 0.070 92.925 ;
    RECT 0 92.995 0.070 93.765 ;
    RECT 0 93.835 0.070 94.605 ;
    RECT 0 94.675 0.070 95.445 ;
    RECT 0 95.515 0.070 96.285 ;
    RECT 0 96.355 0.070 97.125 ;
    RECT 0 97.195 0.070 97.965 ;
    RECT 0 98.035 0.070 98.805 ;
    RECT 0 98.875 0.070 99.645 ;
    RECT 0 99.715 0.070 100.485 ;
    RECT 0 100.555 0.070 101.325 ;
    RECT 0 101.395 0.070 102.165 ;
    RECT 0 102.235 0.070 103.005 ;
    RECT 0 103.075 0.070 103.845 ;
    RECT 0 103.915 0.070 104.685 ;
    RECT 0 104.755 0.070 105.525 ;
    RECT 0 105.595 0.070 106.365 ;
    RECT 0 106.435 0.070 107.205 ;
    RECT 0 107.275 0.070 108.045 ;
    RECT 0 108.115 0.070 108.885 ;
    RECT 0 108.955 0.070 109.725 ;
    RECT 0 109.795 0.070 110.565 ;
    RECT 0 110.635 0.070 111.405 ;
    RECT 0 111.475 0.070 112.245 ;
    RECT 0 112.315 0.070 113.085 ;
    RECT 0 113.155 0.070 113.925 ;
    RECT 0 113.995 0.070 114.765 ;
    RECT 0 114.835 0.070 115.605 ;
    RECT 0 115.675 0.070 116.445 ;
    RECT 0 116.515 0.070 117.285 ;
    RECT 0 117.355 0.070 118.125 ;
    RECT 0 118.195 0.070 118.965 ;
    RECT 0 119.035 0.070 119.805 ;
    RECT 0 119.875 0.070 120.645 ;
    RECT 0 120.715 0.070 121.485 ;
    RECT 0 121.555 0.070 122.325 ;
    RECT 0 122.395 0.070 123.165 ;
    RECT 0 123.235 0.070 124.005 ;
    RECT 0 124.075 0.070 124.845 ;
    RECT 0 124.915 0.070 125.685 ;
    RECT 0 125.755 0.070 126.525 ;
    RECT 0 126.595 0.070 127.365 ;
    RECT 0 127.435 0.070 128.205 ;
    RECT 0 128.275 0.070 129.045 ;
    RECT 0 129.115 0.070 129.885 ;
    RECT 0 129.955 0.070 130.725 ;
    RECT 0 130.795 0.070 131.565 ;
    RECT 0 131.635 0.070 132.405 ;
    RECT 0 132.475 0.070 133.245 ;
    RECT 0 133.315 0.070 134.085 ;
    RECT 0 134.155 0.070 134.925 ;
    RECT 0 134.995 0.070 135.765 ;
    RECT 0 135.835 0.070 136.605 ;
    RECT 0 136.675 0.070 137.445 ;
    RECT 0 137.515 0.070 138.285 ;
    RECT 0 138.355 0.070 139.125 ;
    RECT 0 139.195 0.070 139.965 ;
    RECT 0 140.035 0.070 140.805 ;
    RECT 0 140.875 0.070 141.645 ;
    RECT 0 141.715 0.070 142.485 ;
    RECT 0 142.555 0.070 143.325 ;
    RECT 0 143.395 0.070 144.165 ;
    RECT 0 144.235 0.070 145.005 ;
    RECT 0 145.075 0.070 145.845 ;
    RECT 0 145.915 0.070 146.685 ;
    RECT 0 146.755 0.070 147.525 ;
    RECT 0 147.595 0.070 148.365 ;
    RECT 0 148.435 0.070 149.205 ;
    RECT 0 149.275 0.070 150.045 ;
    RECT 0 150.115 0.070 150.885 ;
    RECT 0 150.955 0.070 151.725 ;
    RECT 0 151.795 0.070 152.565 ;
    RECT 0 152.635 0.070 153.405 ;
    RECT 0 153.475 0.070 154.245 ;
    RECT 0 154.315 0.070 155.085 ;
    RECT 0 155.155 0.070 155.925 ;
    RECT 0 155.995 0.070 156.765 ;
    RECT 0 156.835 0.070 157.605 ;
    RECT 0 157.675 0.070 158.445 ;
    RECT 0 158.515 0.070 159.285 ;
    RECT 0 159.355 0.070 160.125 ;
    RECT 0 160.195 0.070 160.965 ;
    RECT 0 161.035 0.070 161.805 ;
    RECT 0 161.875 0.070 162.645 ;
    RECT 0 162.715 0.070 163.485 ;
    RECT 0 163.555 0.070 164.325 ;
    RECT 0 164.395 0.070 165.165 ;
    RECT 0 165.235 0.070 166.005 ;
    RECT 0 166.075 0.070 166.845 ;
    RECT 0 166.915 0.070 167.685 ;
    RECT 0 167.755 0.070 168.525 ;
    RECT 0 168.595 0.070 169.365 ;
    RECT 0 169.435 0.070 170.205 ;
    RECT 0 170.275 0.070 171.045 ;
    RECT 0 171.115 0.070 171.885 ;
    RECT 0 171.955 0.070 172.725 ;
    RECT 0 172.795 0.070 173.565 ;
    RECT 0 173.635 0.070 174.405 ;
    RECT 0 174.475 0.070 175.245 ;
    RECT 0 175.315 0.070 176.085 ;
    RECT 0 176.155 0.070 176.925 ;
    RECT 0 176.995 0.070 177.765 ;
    RECT 0 177.835 0.070 178.605 ;
    RECT 0 178.675 0.070 179.445 ;
    RECT 0 179.515 0.070 180.285 ;
    RECT 0 180.355 0.070 181.125 ;
    RECT 0 181.195 0.070 181.965 ;
    RECT 0 182.035 0.070 182.805 ;
    RECT 0 182.875 0.070 183.645 ;
    RECT 0 183.715 0.070 184.485 ;
    RECT 0 184.555 0.070 185.325 ;
    RECT 0 185.395 0.070 186.165 ;
    RECT 0 186.235 0.070 187.005 ;
    RECT 0 187.075 0.070 187.845 ;
    RECT 0 187.915 0.070 188.685 ;
    RECT 0 188.755 0.070 189.525 ;
    RECT 0 189.595 0.070 190.365 ;
    RECT 0 190.435 0.070 191.205 ;
    RECT 0 191.275 0.070 192.045 ;
    RECT 0 192.115 0.070 192.885 ;
    RECT 0 192.955 0.070 193.725 ;
    RECT 0 193.795 0.070 194.565 ;
    RECT 0 194.635 0.070 195.405 ;
    RECT 0 195.475 0.070 196.245 ;
    RECT 0 196.315 0.070 197.085 ;
    RECT 0 197.155 0.070 197.925 ;
    RECT 0 197.995 0.070 198.765 ;
    RECT 0 198.835 0.070 199.605 ;
    RECT 0 199.675 0.070 200.445 ;
    RECT 0 200.515 0.070 201.285 ;
    RECT 0 201.355 0.070 202.125 ;
    RECT 0 202.195 0.070 202.965 ;
    RECT 0 203.035 0.070 203.805 ;
    RECT 0 203.875 0.070 204.645 ;
    RECT 0 204.715 0.070 205.485 ;
    RECT 0 205.555 0.070 206.325 ;
    RECT 0 206.395 0.070 207.165 ;
    RECT 0 207.235 0.070 208.005 ;
    RECT 0 208.075 0.070 208.845 ;
    RECT 0 208.915 0.070 209.685 ;
    RECT 0 209.755 0.070 210.525 ;
    RECT 0 210.595 0.070 211.365 ;
    RECT 0 211.435 0.070 212.205 ;
    RECT 0 212.275 0.070 213.045 ;
    RECT 0 213.115 0.070 213.885 ;
    RECT 0 213.955 0.070 214.725 ;
    RECT 0 214.795 0.070 215.565 ;
    RECT 0 215.635 0.070 234.745 ;
    RECT 0 234.815 0.070 235.585 ;
    RECT 0 235.655 0.070 236.425 ;
    RECT 0 236.495 0.070 237.265 ;
    RECT 0 237.335 0.070 238.105 ;
    RECT 0 238.175 0.070 238.945 ;
    RECT 0 239.015 0.070 239.785 ;
    RECT 0 239.855 0.070 240.625 ;
    RECT 0 240.695 0.070 241.465 ;
    RECT 0 241.535 0.070 242.305 ;
    RECT 0 242.375 0.070 243.145 ;
    RECT 0 243.215 0.070 243.985 ;
    RECT 0 244.055 0.070 244.825 ;
    RECT 0 244.895 0.070 245.665 ;
    RECT 0 245.735 0.070 246.505 ;
    RECT 0 246.575 0.070 247.345 ;
    RECT 0 247.415 0.070 248.185 ;
    RECT 0 248.255 0.070 249.025 ;
    RECT 0 249.095 0.070 249.865 ;
    RECT 0 249.935 0.070 250.705 ;
    RECT 0 250.775 0.070 251.545 ;
    RECT 0 251.615 0.070 252.385 ;
    RECT 0 252.455 0.070 253.225 ;
    RECT 0 253.295 0.070 254.065 ;
    RECT 0 254.135 0.070 254.905 ;
    RECT 0 254.975 0.070 255.745 ;
    RECT 0 255.815 0.070 256.585 ;
    RECT 0 256.655 0.070 257.425 ;
    RECT 0 257.495 0.070 258.265 ;
    RECT 0 258.335 0.070 259.105 ;
    RECT 0 259.175 0.070 259.945 ;
    RECT 0 260.015 0.070 260.785 ;
    RECT 0 260.855 0.070 261.625 ;
    RECT 0 261.695 0.070 262.465 ;
    RECT 0 262.535 0.070 263.305 ;
    RECT 0 263.375 0.070 264.145 ;
    RECT 0 264.215 0.070 264.985 ;
    RECT 0 265.055 0.070 265.825 ;
    RECT 0 265.895 0.070 266.665 ;
    RECT 0 266.735 0.070 267.505 ;
    RECT 0 267.575 0.070 268.345 ;
    RECT 0 268.415 0.070 269.185 ;
    RECT 0 269.255 0.070 270.025 ;
    RECT 0 270.095 0.070 270.865 ;
    RECT 0 270.935 0.070 271.705 ;
    RECT 0 271.775 0.070 272.545 ;
    RECT 0 272.615 0.070 273.385 ;
    RECT 0 273.455 0.070 274.225 ;
    RECT 0 274.295 0.070 275.065 ;
    RECT 0 275.135 0.070 275.905 ;
    RECT 0 275.975 0.070 276.745 ;
    RECT 0 276.815 0.070 277.585 ;
    RECT 0 277.655 0.070 278.425 ;
    RECT 0 278.495 0.070 279.265 ;
    RECT 0 279.335 0.070 280.105 ;
    RECT 0 280.175 0.070 280.945 ;
    RECT 0 281.015 0.070 281.785 ;
    RECT 0 281.855 0.070 282.625 ;
    RECT 0 282.695 0.070 283.465 ;
    RECT 0 283.535 0.070 284.305 ;
    RECT 0 284.375 0.070 285.145 ;
    RECT 0 285.215 0.070 285.985 ;
    RECT 0 286.055 0.070 286.825 ;
    RECT 0 286.895 0.070 287.665 ;
    RECT 0 287.735 0.070 288.505 ;
    RECT 0 288.575 0.070 289.345 ;
    RECT 0 289.415 0.070 290.185 ;
    RECT 0 290.255 0.070 291.025 ;
    RECT 0 291.095 0.070 291.865 ;
    RECT 0 291.935 0.070 292.705 ;
    RECT 0 292.775 0.070 293.545 ;
    RECT 0 293.615 0.070 294.385 ;
    RECT 0 294.455 0.070 295.225 ;
    RECT 0 295.295 0.070 296.065 ;
    RECT 0 296.135 0.070 296.905 ;
    RECT 0 296.975 0.070 297.745 ;
    RECT 0 297.815 0.070 298.585 ;
    RECT 0 298.655 0.070 299.425 ;
    RECT 0 299.495 0.070 300.265 ;
    RECT 0 300.335 0.070 301.105 ;
    RECT 0 301.175 0.070 301.945 ;
    RECT 0 302.015 0.070 302.785 ;
    RECT 0 302.855 0.070 303.625 ;
    RECT 0 303.695 0.070 304.465 ;
    RECT 0 304.535 0.070 305.305 ;
    RECT 0 305.375 0.070 306.145 ;
    RECT 0 306.215 0.070 306.985 ;
    RECT 0 307.055 0.070 307.825 ;
    RECT 0 307.895 0.070 308.665 ;
    RECT 0 308.735 0.070 309.505 ;
    RECT 0 309.575 0.070 310.345 ;
    RECT 0 310.415 0.070 311.185 ;
    RECT 0 311.255 0.070 312.025 ;
    RECT 0 312.095 0.070 312.865 ;
    RECT 0 312.935 0.070 313.705 ;
    RECT 0 313.775 0.070 314.545 ;
    RECT 0 314.615 0.070 315.385 ;
    RECT 0 315.455 0.070 316.225 ;
    RECT 0 316.295 0.070 317.065 ;
    RECT 0 317.135 0.070 317.905 ;
    RECT 0 317.975 0.070 318.745 ;
    RECT 0 318.815 0.070 319.585 ;
    RECT 0 319.655 0.070 320.425 ;
    RECT 0 320.495 0.070 321.265 ;
    RECT 0 321.335 0.070 322.105 ;
    RECT 0 322.175 0.070 322.945 ;
    RECT 0 323.015 0.070 323.785 ;
    RECT 0 323.855 0.070 324.625 ;
    RECT 0 324.695 0.070 325.465 ;
    RECT 0 325.535 0.070 326.305 ;
    RECT 0 326.375 0.070 327.145 ;
    RECT 0 327.215 0.070 327.985 ;
    RECT 0 328.055 0.070 328.825 ;
    RECT 0 328.895 0.070 329.665 ;
    RECT 0 329.735 0.070 330.505 ;
    RECT 0 330.575 0.070 331.345 ;
    RECT 0 331.415 0.070 332.185 ;
    RECT 0 332.255 0.070 333.025 ;
    RECT 0 333.095 0.070 333.865 ;
    RECT 0 333.935 0.070 334.705 ;
    RECT 0 334.775 0.070 335.545 ;
    RECT 0 335.615 0.070 336.385 ;
    RECT 0 336.455 0.070 337.225 ;
    RECT 0 337.295 0.070 338.065 ;
    RECT 0 338.135 0.070 338.905 ;
    RECT 0 338.975 0.070 339.745 ;
    RECT 0 339.815 0.070 340.585 ;
    RECT 0 340.655 0.070 341.425 ;
    RECT 0 341.495 0.070 342.265 ;
    RECT 0 342.335 0.070 343.105 ;
    RECT 0 343.175 0.070 343.945 ;
    RECT 0 344.015 0.070 344.785 ;
    RECT 0 344.855 0.070 345.625 ;
    RECT 0 345.695 0.070 346.465 ;
    RECT 0 346.535 0.070 347.305 ;
    RECT 0 347.375 0.070 348.145 ;
    RECT 0 348.215 0.070 348.985 ;
    RECT 0 349.055 0.070 349.825 ;
    RECT 0 349.895 0.070 350.665 ;
    RECT 0 350.735 0.070 351.505 ;
    RECT 0 351.575 0.070 352.345 ;
    RECT 0 352.415 0.070 353.185 ;
    RECT 0 353.255 0.070 354.025 ;
    RECT 0 354.095 0.070 354.865 ;
    RECT 0 354.935 0.070 355.705 ;
    RECT 0 355.775 0.070 356.545 ;
    RECT 0 356.615 0.070 357.385 ;
    RECT 0 357.455 0.070 358.225 ;
    RECT 0 358.295 0.070 359.065 ;
    RECT 0 359.135 0.070 359.905 ;
    RECT 0 359.975 0.070 360.745 ;
    RECT 0 360.815 0.070 361.585 ;
    RECT 0 361.655 0.070 362.425 ;
    RECT 0 362.495 0.070 363.265 ;
    RECT 0 363.335 0.070 364.105 ;
    RECT 0 364.175 0.070 364.945 ;
    RECT 0 365.015 0.070 365.785 ;
    RECT 0 365.855 0.070 366.625 ;
    RECT 0 366.695 0.070 367.465 ;
    RECT 0 367.535 0.070 368.305 ;
    RECT 0 368.375 0.070 369.145 ;
    RECT 0 369.215 0.070 369.985 ;
    RECT 0 370.055 0.070 370.825 ;
    RECT 0 370.895 0.070 371.665 ;
    RECT 0 371.735 0.070 372.505 ;
    RECT 0 372.575 0.070 373.345 ;
    RECT 0 373.415 0.070 374.185 ;
    RECT 0 374.255 0.070 375.025 ;
    RECT 0 375.095 0.070 375.865 ;
    RECT 0 375.935 0.070 376.705 ;
    RECT 0 376.775 0.070 377.545 ;
    RECT 0 377.615 0.070 378.385 ;
    RECT 0 378.455 0.070 379.225 ;
    RECT 0 379.295 0.070 380.065 ;
    RECT 0 380.135 0.070 380.905 ;
    RECT 0 380.975 0.070 381.745 ;
    RECT 0 381.815 0.070 382.585 ;
    RECT 0 382.655 0.070 383.425 ;
    RECT 0 383.495 0.070 384.265 ;
    RECT 0 384.335 0.070 385.105 ;
    RECT 0 385.175 0.070 385.945 ;
    RECT 0 386.015 0.070 386.785 ;
    RECT 0 386.855 0.070 387.625 ;
    RECT 0 387.695 0.070 388.465 ;
    RECT 0 388.535 0.070 389.305 ;
    RECT 0 389.375 0.070 390.145 ;
    RECT 0 390.215 0.070 390.985 ;
    RECT 0 391.055 0.070 391.825 ;
    RECT 0 391.895 0.070 392.665 ;
    RECT 0 392.735 0.070 393.505 ;
    RECT 0 393.575 0.070 394.345 ;
    RECT 0 394.415 0.070 395.185 ;
    RECT 0 395.255 0.070 396.025 ;
    RECT 0 396.095 0.070 396.865 ;
    RECT 0 396.935 0.070 397.705 ;
    RECT 0 397.775 0.070 398.545 ;
    RECT 0 398.615 0.070 399.385 ;
    RECT 0 399.455 0.070 400.225 ;
    RECT 0 400.295 0.070 401.065 ;
    RECT 0 401.135 0.070 401.905 ;
    RECT 0 401.975 0.070 402.745 ;
    RECT 0 402.815 0.070 403.585 ;
    RECT 0 403.655 0.070 404.425 ;
    RECT 0 404.495 0.070 405.265 ;
    RECT 0 405.335 0.070 406.105 ;
    RECT 0 406.175 0.070 406.945 ;
    RECT 0 407.015 0.070 407.785 ;
    RECT 0 407.855 0.070 408.625 ;
    RECT 0 408.695 0.070 409.465 ;
    RECT 0 409.535 0.070 410.305 ;
    RECT 0 410.375 0.070 411.145 ;
    RECT 0 411.215 0.070 411.985 ;
    RECT 0 412.055 0.070 412.825 ;
    RECT 0 412.895 0.070 413.665 ;
    RECT 0 413.735 0.070 414.505 ;
    RECT 0 414.575 0.070 415.345 ;
    RECT 0 415.415 0.070 416.185 ;
    RECT 0 416.255 0.070 417.025 ;
    RECT 0 417.095 0.070 417.865 ;
    RECT 0 417.935 0.070 418.705 ;
    RECT 0 418.775 0.070 419.545 ;
    RECT 0 419.615 0.070 420.385 ;
    RECT 0 420.455 0.070 421.225 ;
    RECT 0 421.295 0.070 422.065 ;
    RECT 0 422.135 0.070 422.905 ;
    RECT 0 422.975 0.070 423.745 ;
    RECT 0 423.815 0.070 424.585 ;
    RECT 0 424.655 0.070 425.425 ;
    RECT 0 425.495 0.070 426.265 ;
    RECT 0 426.335 0.070 427.105 ;
    RECT 0 427.175 0.070 427.945 ;
    RECT 0 428.015 0.070 428.785 ;
    RECT 0 428.855 0.070 429.625 ;
    RECT 0 429.695 0.070 430.465 ;
    RECT 0 430.535 0.070 431.305 ;
    RECT 0 431.375 0.070 432.145 ;
    RECT 0 432.215 0.070 432.985 ;
    RECT 0 433.055 0.070 433.825 ;
    RECT 0 433.895 0.070 434.665 ;
    RECT 0 434.735 0.070 435.505 ;
    RECT 0 435.575 0.070 436.345 ;
    RECT 0 436.415 0.070 437.185 ;
    RECT 0 437.255 0.070 438.025 ;
    RECT 0 438.095 0.070 438.865 ;
    RECT 0 438.935 0.070 439.705 ;
    RECT 0 439.775 0.070 440.545 ;
    RECT 0 440.615 0.070 441.385 ;
    RECT 0 441.455 0.070 442.225 ;
    RECT 0 442.295 0.070 443.065 ;
    RECT 0 443.135 0.070 443.905 ;
    RECT 0 443.975 0.070 444.745 ;
    RECT 0 444.815 0.070 445.585 ;
    RECT 0 445.655 0.070 446.425 ;
    RECT 0 446.495 0.070 447.265 ;
    RECT 0 447.335 0.070 448.105 ;
    RECT 0 448.175 0.070 448.945 ;
    RECT 0 449.015 0.070 468.125 ;
    RECT 0 468.195 0.070 468.965 ;
    RECT 0 469.035 0.070 469.805 ;
    RECT 0 469.875 0.070 470.645 ;
    RECT 0 470.715 0.070 471.485 ;
    RECT 0 471.555 0.070 472.325 ;
    RECT 0 472.395 0.070 473.165 ;
    RECT 0 473.235 0.070 474.005 ;
    RECT 0 474.075 0.070 474.845 ;
    RECT 0 474.915 0.070 475.685 ;
    RECT 0 475.755 0.070 476.525 ;
    RECT 0 476.595 0.070 477.365 ;
    RECT 0 477.435 0.070 478.205 ;
    RECT 0 478.275 0.070 479.045 ;
    RECT 0 479.115 0.070 479.885 ;
    RECT 0 479.955 0.070 480.725 ;
    RECT 0 480.795 0.070 481.565 ;
    RECT 0 481.635 0.070 482.405 ;
    RECT 0 482.475 0.070 483.245 ;
    RECT 0 483.315 0.070 484.085 ;
    RECT 0 484.155 0.070 484.925 ;
    RECT 0 484.995 0.070 485.765 ;
    RECT 0 485.835 0.070 486.605 ;
    RECT 0 486.675 0.070 487.445 ;
    RECT 0 487.515 0.070 488.285 ;
    RECT 0 488.355 0.070 489.125 ;
    RECT 0 489.195 0.070 489.965 ;
    RECT 0 490.035 0.070 490.805 ;
    RECT 0 490.875 0.070 491.645 ;
    RECT 0 491.715 0.070 492.485 ;
    RECT 0 492.555 0.070 493.325 ;
    RECT 0 493.395 0.070 494.165 ;
    RECT 0 494.235 0.070 495.005 ;
    RECT 0 495.075 0.070 495.845 ;
    RECT 0 495.915 0.070 496.685 ;
    RECT 0 496.755 0.070 497.525 ;
    RECT 0 497.595 0.070 498.365 ;
    RECT 0 498.435 0.070 499.205 ;
    RECT 0 499.275 0.070 500.045 ;
    RECT 0 500.115 0.070 500.885 ;
    RECT 0 500.955 0.070 501.725 ;
    RECT 0 501.795 0.070 502.565 ;
    RECT 0 502.635 0.070 503.405 ;
    RECT 0 503.475 0.070 504.245 ;
    RECT 0 504.315 0.070 505.085 ;
    RECT 0 505.155 0.070 505.925 ;
    RECT 0 505.995 0.070 506.765 ;
    RECT 0 506.835 0.070 507.605 ;
    RECT 0 507.675 0.070 508.445 ;
    RECT 0 508.515 0.070 509.285 ;
    RECT 0 509.355 0.070 510.125 ;
    RECT 0 510.195 0.070 510.965 ;
    RECT 0 511.035 0.070 511.805 ;
    RECT 0 511.875 0.070 512.645 ;
    RECT 0 512.715 0.070 513.485 ;
    RECT 0 513.555 0.070 514.325 ;
    RECT 0 514.395 0.070 515.165 ;
    RECT 0 515.235 0.070 516.005 ;
    RECT 0 516.075 0.070 516.845 ;
    RECT 0 516.915 0.070 517.685 ;
    RECT 0 517.755 0.070 518.525 ;
    RECT 0 518.595 0.070 519.365 ;
    RECT 0 519.435 0.070 520.205 ;
    RECT 0 520.275 0.070 521.045 ;
    RECT 0 521.115 0.070 521.885 ;
    RECT 0 521.955 0.070 522.725 ;
    RECT 0 522.795 0.070 523.565 ;
    RECT 0 523.635 0.070 524.405 ;
    RECT 0 524.475 0.070 525.245 ;
    RECT 0 525.315 0.070 526.085 ;
    RECT 0 526.155 0.070 526.925 ;
    RECT 0 526.995 0.070 527.765 ;
    RECT 0 527.835 0.070 528.605 ;
    RECT 0 528.675 0.070 529.445 ;
    RECT 0 529.515 0.070 530.285 ;
    RECT 0 530.355 0.070 531.125 ;
    RECT 0 531.195 0.070 531.965 ;
    RECT 0 532.035 0.070 532.805 ;
    RECT 0 532.875 0.070 533.645 ;
    RECT 0 533.715 0.070 534.485 ;
    RECT 0 534.555 0.070 535.325 ;
    RECT 0 535.395 0.070 536.165 ;
    RECT 0 536.235 0.070 537.005 ;
    RECT 0 537.075 0.070 537.845 ;
    RECT 0 537.915 0.070 538.685 ;
    RECT 0 538.755 0.070 539.525 ;
    RECT 0 539.595 0.070 540.365 ;
    RECT 0 540.435 0.070 541.205 ;
    RECT 0 541.275 0.070 542.045 ;
    RECT 0 542.115 0.070 542.885 ;
    RECT 0 542.955 0.070 543.725 ;
    RECT 0 543.795 0.070 544.565 ;
    RECT 0 544.635 0.070 545.405 ;
    RECT 0 545.475 0.070 546.245 ;
    RECT 0 546.315 0.070 547.085 ;
    RECT 0 547.155 0.070 547.925 ;
    RECT 0 547.995 0.070 548.765 ;
    RECT 0 548.835 0.070 549.605 ;
    RECT 0 549.675 0.070 550.445 ;
    RECT 0 550.515 0.070 551.285 ;
    RECT 0 551.355 0.070 552.125 ;
    RECT 0 552.195 0.070 552.965 ;
    RECT 0 553.035 0.070 553.805 ;
    RECT 0 553.875 0.070 554.645 ;
    RECT 0 554.715 0.070 555.485 ;
    RECT 0 555.555 0.070 556.325 ;
    RECT 0 556.395 0.070 557.165 ;
    RECT 0 557.235 0.070 558.005 ;
    RECT 0 558.075 0.070 558.845 ;
    RECT 0 558.915 0.070 559.685 ;
    RECT 0 559.755 0.070 560.525 ;
    RECT 0 560.595 0.070 561.365 ;
    RECT 0 561.435 0.070 562.205 ;
    RECT 0 562.275 0.070 563.045 ;
    RECT 0 563.115 0.070 563.885 ;
    RECT 0 563.955 0.070 564.725 ;
    RECT 0 564.795 0.070 565.565 ;
    RECT 0 565.635 0.070 566.405 ;
    RECT 0 566.475 0.070 567.245 ;
    RECT 0 567.315 0.070 568.085 ;
    RECT 0 568.155 0.070 568.925 ;
    RECT 0 568.995 0.070 569.765 ;
    RECT 0 569.835 0.070 570.605 ;
    RECT 0 570.675 0.070 571.445 ;
    RECT 0 571.515 0.070 572.285 ;
    RECT 0 572.355 0.070 573.125 ;
    RECT 0 573.195 0.070 573.965 ;
    RECT 0 574.035 0.070 574.805 ;
    RECT 0 574.875 0.070 575.645 ;
    RECT 0 575.715 0.070 576.485 ;
    RECT 0 576.555 0.070 577.325 ;
    RECT 0 577.395 0.070 578.165 ;
    RECT 0 578.235 0.070 579.005 ;
    RECT 0 579.075 0.070 579.845 ;
    RECT 0 579.915 0.070 580.685 ;
    RECT 0 580.755 0.070 581.525 ;
    RECT 0 581.595 0.070 582.365 ;
    RECT 0 582.435 0.070 583.205 ;
    RECT 0 583.275 0.070 584.045 ;
    RECT 0 584.115 0.070 584.885 ;
    RECT 0 584.955 0.070 585.725 ;
    RECT 0 585.795 0.070 586.565 ;
    RECT 0 586.635 0.070 587.405 ;
    RECT 0 587.475 0.070 588.245 ;
    RECT 0 588.315 0.070 589.085 ;
    RECT 0 589.155 0.070 589.925 ;
    RECT 0 589.995 0.070 590.765 ;
    RECT 0 590.835 0.070 591.605 ;
    RECT 0 591.675 0.070 592.445 ;
    RECT 0 592.515 0.070 593.285 ;
    RECT 0 593.355 0.070 594.125 ;
    RECT 0 594.195 0.070 594.965 ;
    RECT 0 595.035 0.070 595.805 ;
    RECT 0 595.875 0.070 596.645 ;
    RECT 0 596.715 0.070 597.485 ;
    RECT 0 597.555 0.070 598.325 ;
    RECT 0 598.395 0.070 599.165 ;
    RECT 0 599.235 0.070 600.005 ;
    RECT 0 600.075 0.070 600.845 ;
    RECT 0 600.915 0.070 601.685 ;
    RECT 0 601.755 0.070 602.525 ;
    RECT 0 602.595 0.070 603.365 ;
    RECT 0 603.435 0.070 604.205 ;
    RECT 0 604.275 0.070 605.045 ;
    RECT 0 605.115 0.070 605.885 ;
    RECT 0 605.955 0.070 606.725 ;
    RECT 0 606.795 0.070 607.565 ;
    RECT 0 607.635 0.070 608.405 ;
    RECT 0 608.475 0.070 609.245 ;
    RECT 0 609.315 0.070 610.085 ;
    RECT 0 610.155 0.070 610.925 ;
    RECT 0 610.995 0.070 611.765 ;
    RECT 0 611.835 0.070 612.605 ;
    RECT 0 612.675 0.070 613.445 ;
    RECT 0 613.515 0.070 614.285 ;
    RECT 0 614.355 0.070 615.125 ;
    RECT 0 615.195 0.070 615.965 ;
    RECT 0 616.035 0.070 616.805 ;
    RECT 0 616.875 0.070 617.645 ;
    RECT 0 617.715 0.070 618.485 ;
    RECT 0 618.555 0.070 619.325 ;
    RECT 0 619.395 0.070 620.165 ;
    RECT 0 620.235 0.070 621.005 ;
    RECT 0 621.075 0.070 621.845 ;
    RECT 0 621.915 0.070 622.685 ;
    RECT 0 622.755 0.070 623.525 ;
    RECT 0 623.595 0.070 624.365 ;
    RECT 0 624.435 0.070 625.205 ;
    RECT 0 625.275 0.070 626.045 ;
    RECT 0 626.115 0.070 626.885 ;
    RECT 0 626.955 0.070 627.725 ;
    RECT 0 627.795 0.070 628.565 ;
    RECT 0 628.635 0.070 629.405 ;
    RECT 0 629.475 0.070 630.245 ;
    RECT 0 630.315 0.070 631.085 ;
    RECT 0 631.155 0.070 631.925 ;
    RECT 0 631.995 0.070 632.765 ;
    RECT 0 632.835 0.070 633.605 ;
    RECT 0 633.675 0.070 634.445 ;
    RECT 0 634.515 0.070 635.285 ;
    RECT 0 635.355 0.070 636.125 ;
    RECT 0 636.195 0.070 636.965 ;
    RECT 0 637.035 0.070 637.805 ;
    RECT 0 637.875 0.070 638.645 ;
    RECT 0 638.715 0.070 639.485 ;
    RECT 0 639.555 0.070 640.325 ;
    RECT 0 640.395 0.070 641.165 ;
    RECT 0 641.235 0.070 642.005 ;
    RECT 0 642.075 0.070 642.845 ;
    RECT 0 642.915 0.070 643.685 ;
    RECT 0 643.755 0.070 644.525 ;
    RECT 0 644.595 0.070 645.365 ;
    RECT 0 645.435 0.070 646.205 ;
    RECT 0 646.275 0.070 647.045 ;
    RECT 0 647.115 0.070 647.885 ;
    RECT 0 647.955 0.070 648.725 ;
    RECT 0 648.795 0.070 649.565 ;
    RECT 0 649.635 0.070 650.405 ;
    RECT 0 650.475 0.070 651.245 ;
    RECT 0 651.315 0.070 652.085 ;
    RECT 0 652.155 0.070 652.925 ;
    RECT 0 652.995 0.070 653.765 ;
    RECT 0 653.835 0.070 654.605 ;
    RECT 0 654.675 0.070 655.445 ;
    RECT 0 655.515 0.070 656.285 ;
    RECT 0 656.355 0.070 657.125 ;
    RECT 0 657.195 0.070 657.965 ;
    RECT 0 658.035 0.070 658.805 ;
    RECT 0 658.875 0.070 659.645 ;
    RECT 0 659.715 0.070 660.485 ;
    RECT 0 660.555 0.070 661.325 ;
    RECT 0 661.395 0.070 662.165 ;
    RECT 0 662.235 0.070 663.005 ;
    RECT 0 663.075 0.070 663.845 ;
    RECT 0 663.915 0.070 664.685 ;
    RECT 0 664.755 0.070 665.525 ;
    RECT 0 665.595 0.070 666.365 ;
    RECT 0 666.435 0.070 667.205 ;
    RECT 0 667.275 0.070 668.045 ;
    RECT 0 668.115 0.070 668.885 ;
    RECT 0 668.955 0.070 669.725 ;
    RECT 0 669.795 0.070 670.565 ;
    RECT 0 670.635 0.070 671.405 ;
    RECT 0 671.475 0.070 672.245 ;
    RECT 0 672.315 0.070 673.085 ;
    RECT 0 673.155 0.070 673.925 ;
    RECT 0 673.995 0.070 674.765 ;
    RECT 0 674.835 0.070 675.605 ;
    RECT 0 675.675 0.070 676.445 ;
    RECT 0 676.515 0.070 677.285 ;
    RECT 0 677.355 0.070 678.125 ;
    RECT 0 678.195 0.070 678.965 ;
    RECT 0 679.035 0.070 679.805 ;
    RECT 0 679.875 0.070 680.645 ;
    RECT 0 680.715 0.070 681.485 ;
    RECT 0 681.555 0.070 682.325 ;
    RECT 0 682.395 0.070 701.505 ;
    RECT 0 701.575 0.070 702.345 ;
    RECT 0 702.415 0.070 703.185 ;
    RECT 0 703.255 0.070 704.025 ;
    RECT 0 704.095 0.070 704.865 ;
    RECT 0 704.935 0.070 705.705 ;
    RECT 0 705.775 0.070 706.545 ;
    RECT 0 706.615 0.070 707.385 ;
    RECT 0 707.455 0.070 708.225 ;
    RECT 0 708.295 0.070 709.065 ;
    RECT 0 709.135 0.070 709.905 ;
    RECT 0 709.975 0.070 710.745 ;
    RECT 0 710.815 0.070 729.925 ;
    RECT 0 729.995 0.070 730.765 ;
    RECT 0 730.835 0.070 731.605 ;
    RECT 0 731.675 0.070 737.800 ;
    LAYER metal4 ;
    RECT 0 0 1631.530 1.400 ;
    RECT 0 736.400 1631.530 737.800 ;
    RECT 0.000 1.400 1.260 736.400 ;
    RECT 1.540 1.400 2.380 736.400 ;
    RECT 2.660 1.400 3.500 736.400 ;
    RECT 3.780 1.400 4.620 736.400 ;
    RECT 4.900 1.400 5.740 736.400 ;
    RECT 6.020 1.400 6.860 736.400 ;
    RECT 7.140 1.400 7.980 736.400 ;
    RECT 8.260 1.400 9.100 736.400 ;
    RECT 9.380 1.400 10.220 736.400 ;
    RECT 10.500 1.400 11.340 736.400 ;
    RECT 11.620 1.400 12.460 736.400 ;
    RECT 12.740 1.400 13.580 736.400 ;
    RECT 13.860 1.400 14.700 736.400 ;
    RECT 14.980 1.400 15.820 736.400 ;
    RECT 16.100 1.400 16.940 736.400 ;
    RECT 17.220 1.400 18.060 736.400 ;
    RECT 18.340 1.400 19.180 736.400 ;
    RECT 19.460 1.400 20.300 736.400 ;
    RECT 20.580 1.400 21.420 736.400 ;
    RECT 21.700 1.400 22.540 736.400 ;
    RECT 22.820 1.400 23.660 736.400 ;
    RECT 23.940 1.400 24.780 736.400 ;
    RECT 25.060 1.400 25.900 736.400 ;
    RECT 26.180 1.400 27.020 736.400 ;
    RECT 27.300 1.400 28.140 736.400 ;
    RECT 28.420 1.400 29.260 736.400 ;
    RECT 29.540 1.400 30.380 736.400 ;
    RECT 30.660 1.400 31.500 736.400 ;
    RECT 31.780 1.400 32.620 736.400 ;
    RECT 32.900 1.400 33.740 736.400 ;
    RECT 34.020 1.400 34.860 736.400 ;
    RECT 35.140 1.400 35.980 736.400 ;
    RECT 36.260 1.400 37.100 736.400 ;
    RECT 37.380 1.400 38.220 736.400 ;
    RECT 38.500 1.400 39.340 736.400 ;
    RECT 39.620 1.400 40.460 736.400 ;
    RECT 40.740 1.400 41.580 736.400 ;
    RECT 41.860 1.400 42.700 736.400 ;
    RECT 42.980 1.400 43.820 736.400 ;
    RECT 44.100 1.400 44.940 736.400 ;
    RECT 45.220 1.400 46.060 736.400 ;
    RECT 46.340 1.400 47.180 736.400 ;
    RECT 47.460 1.400 48.300 736.400 ;
    RECT 48.580 1.400 49.420 736.400 ;
    RECT 49.700 1.400 50.540 736.400 ;
    RECT 50.820 1.400 51.660 736.400 ;
    RECT 51.940 1.400 52.780 736.400 ;
    RECT 53.060 1.400 53.900 736.400 ;
    RECT 54.180 1.400 55.020 736.400 ;
    RECT 55.300 1.400 56.140 736.400 ;
    RECT 56.420 1.400 57.260 736.400 ;
    RECT 57.540 1.400 58.380 736.400 ;
    RECT 58.660 1.400 59.500 736.400 ;
    RECT 59.780 1.400 60.620 736.400 ;
    RECT 60.900 1.400 61.740 736.400 ;
    RECT 62.020 1.400 62.860 736.400 ;
    RECT 63.140 1.400 63.980 736.400 ;
    RECT 64.260 1.400 65.100 736.400 ;
    RECT 65.380 1.400 66.220 736.400 ;
    RECT 66.500 1.400 67.340 736.400 ;
    RECT 67.620 1.400 68.460 736.400 ;
    RECT 68.740 1.400 69.580 736.400 ;
    RECT 69.860 1.400 70.700 736.400 ;
    RECT 70.980 1.400 71.820 736.400 ;
    RECT 72.100 1.400 72.940 736.400 ;
    RECT 73.220 1.400 74.060 736.400 ;
    RECT 74.340 1.400 75.180 736.400 ;
    RECT 75.460 1.400 76.300 736.400 ;
    RECT 76.580 1.400 77.420 736.400 ;
    RECT 77.700 1.400 78.540 736.400 ;
    RECT 78.820 1.400 79.660 736.400 ;
    RECT 79.940 1.400 80.780 736.400 ;
    RECT 81.060 1.400 81.900 736.400 ;
    RECT 82.180 1.400 83.020 736.400 ;
    RECT 83.300 1.400 84.140 736.400 ;
    RECT 84.420 1.400 85.260 736.400 ;
    RECT 85.540 1.400 86.380 736.400 ;
    RECT 86.660 1.400 87.500 736.400 ;
    RECT 87.780 1.400 88.620 736.400 ;
    RECT 88.900 1.400 89.740 736.400 ;
    RECT 90.020 1.400 90.860 736.400 ;
    RECT 91.140 1.400 91.980 736.400 ;
    RECT 92.260 1.400 93.100 736.400 ;
    RECT 93.380 1.400 94.220 736.400 ;
    RECT 94.500 1.400 95.340 736.400 ;
    RECT 95.620 1.400 96.460 736.400 ;
    RECT 96.740 1.400 97.580 736.400 ;
    RECT 97.860 1.400 98.700 736.400 ;
    RECT 98.980 1.400 99.820 736.400 ;
    RECT 100.100 1.400 100.940 736.400 ;
    RECT 101.220 1.400 102.060 736.400 ;
    RECT 102.340 1.400 103.180 736.400 ;
    RECT 103.460 1.400 104.300 736.400 ;
    RECT 104.580 1.400 105.420 736.400 ;
    RECT 105.700 1.400 106.540 736.400 ;
    RECT 106.820 1.400 107.660 736.400 ;
    RECT 107.940 1.400 108.780 736.400 ;
    RECT 109.060 1.400 109.900 736.400 ;
    RECT 110.180 1.400 111.020 736.400 ;
    RECT 111.300 1.400 112.140 736.400 ;
    RECT 112.420 1.400 113.260 736.400 ;
    RECT 113.540 1.400 114.380 736.400 ;
    RECT 114.660 1.400 115.500 736.400 ;
    RECT 115.780 1.400 116.620 736.400 ;
    RECT 116.900 1.400 117.740 736.400 ;
    RECT 118.020 1.400 118.860 736.400 ;
    RECT 119.140 1.400 119.980 736.400 ;
    RECT 120.260 1.400 121.100 736.400 ;
    RECT 121.380 1.400 122.220 736.400 ;
    RECT 122.500 1.400 123.340 736.400 ;
    RECT 123.620 1.400 124.460 736.400 ;
    RECT 124.740 1.400 125.580 736.400 ;
    RECT 125.860 1.400 126.700 736.400 ;
    RECT 126.980 1.400 127.820 736.400 ;
    RECT 128.100 1.400 128.940 736.400 ;
    RECT 129.220 1.400 130.060 736.400 ;
    RECT 130.340 1.400 131.180 736.400 ;
    RECT 131.460 1.400 132.300 736.400 ;
    RECT 132.580 1.400 133.420 736.400 ;
    RECT 133.700 1.400 134.540 736.400 ;
    RECT 134.820 1.400 135.660 736.400 ;
    RECT 135.940 1.400 136.780 736.400 ;
    RECT 137.060 1.400 137.900 736.400 ;
    RECT 138.180 1.400 139.020 736.400 ;
    RECT 139.300 1.400 140.140 736.400 ;
    RECT 140.420 1.400 141.260 736.400 ;
    RECT 141.540 1.400 142.380 736.400 ;
    RECT 142.660 1.400 143.500 736.400 ;
    RECT 143.780 1.400 144.620 736.400 ;
    RECT 144.900 1.400 145.740 736.400 ;
    RECT 146.020 1.400 146.860 736.400 ;
    RECT 147.140 1.400 147.980 736.400 ;
    RECT 148.260 1.400 149.100 736.400 ;
    RECT 149.380 1.400 150.220 736.400 ;
    RECT 150.500 1.400 151.340 736.400 ;
    RECT 151.620 1.400 152.460 736.400 ;
    RECT 152.740 1.400 153.580 736.400 ;
    RECT 153.860 1.400 154.700 736.400 ;
    RECT 154.980 1.400 155.820 736.400 ;
    RECT 156.100 1.400 156.940 736.400 ;
    RECT 157.220 1.400 158.060 736.400 ;
    RECT 158.340 1.400 159.180 736.400 ;
    RECT 159.460 1.400 160.300 736.400 ;
    RECT 160.580 1.400 161.420 736.400 ;
    RECT 161.700 1.400 162.540 736.400 ;
    RECT 162.820 1.400 163.660 736.400 ;
    RECT 163.940 1.400 164.780 736.400 ;
    RECT 165.060 1.400 165.900 736.400 ;
    RECT 166.180 1.400 167.020 736.400 ;
    RECT 167.300 1.400 168.140 736.400 ;
    RECT 168.420 1.400 169.260 736.400 ;
    RECT 169.540 1.400 170.380 736.400 ;
    RECT 170.660 1.400 171.500 736.400 ;
    RECT 171.780 1.400 172.620 736.400 ;
    RECT 172.900 1.400 173.740 736.400 ;
    RECT 174.020 1.400 174.860 736.400 ;
    RECT 175.140 1.400 175.980 736.400 ;
    RECT 176.260 1.400 177.100 736.400 ;
    RECT 177.380 1.400 178.220 736.400 ;
    RECT 178.500 1.400 179.340 736.400 ;
    RECT 179.620 1.400 180.460 736.400 ;
    RECT 180.740 1.400 181.580 736.400 ;
    RECT 181.860 1.400 182.700 736.400 ;
    RECT 182.980 1.400 183.820 736.400 ;
    RECT 184.100 1.400 184.940 736.400 ;
    RECT 185.220 1.400 186.060 736.400 ;
    RECT 186.340 1.400 187.180 736.400 ;
    RECT 187.460 1.400 188.300 736.400 ;
    RECT 188.580 1.400 189.420 736.400 ;
    RECT 189.700 1.400 190.540 736.400 ;
    RECT 190.820 1.400 191.660 736.400 ;
    RECT 191.940 1.400 192.780 736.400 ;
    RECT 193.060 1.400 193.900 736.400 ;
    RECT 194.180 1.400 195.020 736.400 ;
    RECT 195.300 1.400 196.140 736.400 ;
    RECT 196.420 1.400 197.260 736.400 ;
    RECT 197.540 1.400 198.380 736.400 ;
    RECT 198.660 1.400 199.500 736.400 ;
    RECT 199.780 1.400 200.620 736.400 ;
    RECT 200.900 1.400 201.740 736.400 ;
    RECT 202.020 1.400 202.860 736.400 ;
    RECT 203.140 1.400 203.980 736.400 ;
    RECT 204.260 1.400 205.100 736.400 ;
    RECT 205.380 1.400 206.220 736.400 ;
    RECT 206.500 1.400 207.340 736.400 ;
    RECT 207.620 1.400 208.460 736.400 ;
    RECT 208.740 1.400 209.580 736.400 ;
    RECT 209.860 1.400 210.700 736.400 ;
    RECT 210.980 1.400 211.820 736.400 ;
    RECT 212.100 1.400 212.940 736.400 ;
    RECT 213.220 1.400 214.060 736.400 ;
    RECT 214.340 1.400 215.180 736.400 ;
    RECT 215.460 1.400 216.300 736.400 ;
    RECT 216.580 1.400 217.420 736.400 ;
    RECT 217.700 1.400 218.540 736.400 ;
    RECT 218.820 1.400 219.660 736.400 ;
    RECT 219.940 1.400 220.780 736.400 ;
    RECT 221.060 1.400 221.900 736.400 ;
    RECT 222.180 1.400 223.020 736.400 ;
    RECT 223.300 1.400 224.140 736.400 ;
    RECT 224.420 1.400 225.260 736.400 ;
    RECT 225.540 1.400 226.380 736.400 ;
    RECT 226.660 1.400 227.500 736.400 ;
    RECT 227.780 1.400 228.620 736.400 ;
    RECT 228.900 1.400 229.740 736.400 ;
    RECT 230.020 1.400 230.860 736.400 ;
    RECT 231.140 1.400 231.980 736.400 ;
    RECT 232.260 1.400 233.100 736.400 ;
    RECT 233.380 1.400 234.220 736.400 ;
    RECT 234.500 1.400 235.340 736.400 ;
    RECT 235.620 1.400 236.460 736.400 ;
    RECT 236.740 1.400 237.580 736.400 ;
    RECT 237.860 1.400 238.700 736.400 ;
    RECT 238.980 1.400 239.820 736.400 ;
    RECT 240.100 1.400 240.940 736.400 ;
    RECT 241.220 1.400 242.060 736.400 ;
    RECT 242.340 1.400 243.180 736.400 ;
    RECT 243.460 1.400 244.300 736.400 ;
    RECT 244.580 1.400 245.420 736.400 ;
    RECT 245.700 1.400 246.540 736.400 ;
    RECT 246.820 1.400 247.660 736.400 ;
    RECT 247.940 1.400 248.780 736.400 ;
    RECT 249.060 1.400 249.900 736.400 ;
    RECT 250.180 1.400 251.020 736.400 ;
    RECT 251.300 1.400 252.140 736.400 ;
    RECT 252.420 1.400 253.260 736.400 ;
    RECT 253.540 1.400 254.380 736.400 ;
    RECT 254.660 1.400 255.500 736.400 ;
    RECT 255.780 1.400 256.620 736.400 ;
    RECT 256.900 1.400 257.740 736.400 ;
    RECT 258.020 1.400 258.860 736.400 ;
    RECT 259.140 1.400 259.980 736.400 ;
    RECT 260.260 1.400 261.100 736.400 ;
    RECT 261.380 1.400 262.220 736.400 ;
    RECT 262.500 1.400 263.340 736.400 ;
    RECT 263.620 1.400 264.460 736.400 ;
    RECT 264.740 1.400 265.580 736.400 ;
    RECT 265.860 1.400 266.700 736.400 ;
    RECT 266.980 1.400 267.820 736.400 ;
    RECT 268.100 1.400 268.940 736.400 ;
    RECT 269.220 1.400 270.060 736.400 ;
    RECT 270.340 1.400 271.180 736.400 ;
    RECT 271.460 1.400 272.300 736.400 ;
    RECT 272.580 1.400 273.420 736.400 ;
    RECT 273.700 1.400 274.540 736.400 ;
    RECT 274.820 1.400 275.660 736.400 ;
    RECT 275.940 1.400 276.780 736.400 ;
    RECT 277.060 1.400 277.900 736.400 ;
    RECT 278.180 1.400 279.020 736.400 ;
    RECT 279.300 1.400 280.140 736.400 ;
    RECT 280.420 1.400 281.260 736.400 ;
    RECT 281.540 1.400 282.380 736.400 ;
    RECT 282.660 1.400 283.500 736.400 ;
    RECT 283.780 1.400 284.620 736.400 ;
    RECT 284.900 1.400 285.740 736.400 ;
    RECT 286.020 1.400 286.860 736.400 ;
    RECT 287.140 1.400 287.980 736.400 ;
    RECT 288.260 1.400 289.100 736.400 ;
    RECT 289.380 1.400 290.220 736.400 ;
    RECT 290.500 1.400 291.340 736.400 ;
    RECT 291.620 1.400 292.460 736.400 ;
    RECT 292.740 1.400 293.580 736.400 ;
    RECT 293.860 1.400 294.700 736.400 ;
    RECT 294.980 1.400 295.820 736.400 ;
    RECT 296.100 1.400 296.940 736.400 ;
    RECT 297.220 1.400 298.060 736.400 ;
    RECT 298.340 1.400 299.180 736.400 ;
    RECT 299.460 1.400 300.300 736.400 ;
    RECT 300.580 1.400 301.420 736.400 ;
    RECT 301.700 1.400 302.540 736.400 ;
    RECT 302.820 1.400 303.660 736.400 ;
    RECT 303.940 1.400 304.780 736.400 ;
    RECT 305.060 1.400 305.900 736.400 ;
    RECT 306.180 1.400 307.020 736.400 ;
    RECT 307.300 1.400 308.140 736.400 ;
    RECT 308.420 1.400 309.260 736.400 ;
    RECT 309.540 1.400 310.380 736.400 ;
    RECT 310.660 1.400 311.500 736.400 ;
    RECT 311.780 1.400 312.620 736.400 ;
    RECT 312.900 1.400 313.740 736.400 ;
    RECT 314.020 1.400 314.860 736.400 ;
    RECT 315.140 1.400 315.980 736.400 ;
    RECT 316.260 1.400 317.100 736.400 ;
    RECT 317.380 1.400 318.220 736.400 ;
    RECT 318.500 1.400 319.340 736.400 ;
    RECT 319.620 1.400 320.460 736.400 ;
    RECT 320.740 1.400 321.580 736.400 ;
    RECT 321.860 1.400 322.700 736.400 ;
    RECT 322.980 1.400 323.820 736.400 ;
    RECT 324.100 1.400 324.940 736.400 ;
    RECT 325.220 1.400 326.060 736.400 ;
    RECT 326.340 1.400 327.180 736.400 ;
    RECT 327.460 1.400 328.300 736.400 ;
    RECT 328.580 1.400 329.420 736.400 ;
    RECT 329.700 1.400 330.540 736.400 ;
    RECT 330.820 1.400 331.660 736.400 ;
    RECT 331.940 1.400 332.780 736.400 ;
    RECT 333.060 1.400 333.900 736.400 ;
    RECT 334.180 1.400 335.020 736.400 ;
    RECT 335.300 1.400 336.140 736.400 ;
    RECT 336.420 1.400 337.260 736.400 ;
    RECT 337.540 1.400 338.380 736.400 ;
    RECT 338.660 1.400 339.500 736.400 ;
    RECT 339.780 1.400 340.620 736.400 ;
    RECT 340.900 1.400 341.740 736.400 ;
    RECT 342.020 1.400 342.860 736.400 ;
    RECT 343.140 1.400 343.980 736.400 ;
    RECT 344.260 1.400 345.100 736.400 ;
    RECT 345.380 1.400 346.220 736.400 ;
    RECT 346.500 1.400 347.340 736.400 ;
    RECT 347.620 1.400 348.460 736.400 ;
    RECT 348.740 1.400 349.580 736.400 ;
    RECT 349.860 1.400 350.700 736.400 ;
    RECT 350.980 1.400 351.820 736.400 ;
    RECT 352.100 1.400 352.940 736.400 ;
    RECT 353.220 1.400 354.060 736.400 ;
    RECT 354.340 1.400 355.180 736.400 ;
    RECT 355.460 1.400 356.300 736.400 ;
    RECT 356.580 1.400 357.420 736.400 ;
    RECT 357.700 1.400 358.540 736.400 ;
    RECT 358.820 1.400 359.660 736.400 ;
    RECT 359.940 1.400 360.780 736.400 ;
    RECT 361.060 1.400 361.900 736.400 ;
    RECT 362.180 1.400 363.020 736.400 ;
    RECT 363.300 1.400 364.140 736.400 ;
    RECT 364.420 1.400 365.260 736.400 ;
    RECT 365.540 1.400 366.380 736.400 ;
    RECT 366.660 1.400 367.500 736.400 ;
    RECT 367.780 1.400 368.620 736.400 ;
    RECT 368.900 1.400 369.740 736.400 ;
    RECT 370.020 1.400 370.860 736.400 ;
    RECT 371.140 1.400 371.980 736.400 ;
    RECT 372.260 1.400 373.100 736.400 ;
    RECT 373.380 1.400 374.220 736.400 ;
    RECT 374.500 1.400 375.340 736.400 ;
    RECT 375.620 1.400 376.460 736.400 ;
    RECT 376.740 1.400 377.580 736.400 ;
    RECT 377.860 1.400 378.700 736.400 ;
    RECT 378.980 1.400 379.820 736.400 ;
    RECT 380.100 1.400 380.940 736.400 ;
    RECT 381.220 1.400 382.060 736.400 ;
    RECT 382.340 1.400 383.180 736.400 ;
    RECT 383.460 1.400 384.300 736.400 ;
    RECT 384.580 1.400 385.420 736.400 ;
    RECT 385.700 1.400 386.540 736.400 ;
    RECT 386.820 1.400 387.660 736.400 ;
    RECT 387.940 1.400 388.780 736.400 ;
    RECT 389.060 1.400 389.900 736.400 ;
    RECT 390.180 1.400 391.020 736.400 ;
    RECT 391.300 1.400 392.140 736.400 ;
    RECT 392.420 1.400 393.260 736.400 ;
    RECT 393.540 1.400 394.380 736.400 ;
    RECT 394.660 1.400 395.500 736.400 ;
    RECT 395.780 1.400 396.620 736.400 ;
    RECT 396.900 1.400 397.740 736.400 ;
    RECT 398.020 1.400 398.860 736.400 ;
    RECT 399.140 1.400 399.980 736.400 ;
    RECT 400.260 1.400 401.100 736.400 ;
    RECT 401.380 1.400 402.220 736.400 ;
    RECT 402.500 1.400 403.340 736.400 ;
    RECT 403.620 1.400 404.460 736.400 ;
    RECT 404.740 1.400 405.580 736.400 ;
    RECT 405.860 1.400 406.700 736.400 ;
    RECT 406.980 1.400 407.820 736.400 ;
    RECT 408.100 1.400 408.940 736.400 ;
    RECT 409.220 1.400 410.060 736.400 ;
    RECT 410.340 1.400 411.180 736.400 ;
    RECT 411.460 1.400 412.300 736.400 ;
    RECT 412.580 1.400 413.420 736.400 ;
    RECT 413.700 1.400 414.540 736.400 ;
    RECT 414.820 1.400 415.660 736.400 ;
    RECT 415.940 1.400 416.780 736.400 ;
    RECT 417.060 1.400 417.900 736.400 ;
    RECT 418.180 1.400 419.020 736.400 ;
    RECT 419.300 1.400 420.140 736.400 ;
    RECT 420.420 1.400 421.260 736.400 ;
    RECT 421.540 1.400 422.380 736.400 ;
    RECT 422.660 1.400 423.500 736.400 ;
    RECT 423.780 1.400 424.620 736.400 ;
    RECT 424.900 1.400 425.740 736.400 ;
    RECT 426.020 1.400 426.860 736.400 ;
    RECT 427.140 1.400 427.980 736.400 ;
    RECT 428.260 1.400 429.100 736.400 ;
    RECT 429.380 1.400 430.220 736.400 ;
    RECT 430.500 1.400 431.340 736.400 ;
    RECT 431.620 1.400 432.460 736.400 ;
    RECT 432.740 1.400 433.580 736.400 ;
    RECT 433.860 1.400 434.700 736.400 ;
    RECT 434.980 1.400 435.820 736.400 ;
    RECT 436.100 1.400 436.940 736.400 ;
    RECT 437.220 1.400 438.060 736.400 ;
    RECT 438.340 1.400 439.180 736.400 ;
    RECT 439.460 1.400 440.300 736.400 ;
    RECT 440.580 1.400 441.420 736.400 ;
    RECT 441.700 1.400 442.540 736.400 ;
    RECT 442.820 1.400 443.660 736.400 ;
    RECT 443.940 1.400 444.780 736.400 ;
    RECT 445.060 1.400 445.900 736.400 ;
    RECT 446.180 1.400 447.020 736.400 ;
    RECT 447.300 1.400 448.140 736.400 ;
    RECT 448.420 1.400 449.260 736.400 ;
    RECT 449.540 1.400 450.380 736.400 ;
    RECT 450.660 1.400 451.500 736.400 ;
    RECT 451.780 1.400 452.620 736.400 ;
    RECT 452.900 1.400 453.740 736.400 ;
    RECT 454.020 1.400 454.860 736.400 ;
    RECT 455.140 1.400 455.980 736.400 ;
    RECT 456.260 1.400 457.100 736.400 ;
    RECT 457.380 1.400 458.220 736.400 ;
    RECT 458.500 1.400 459.340 736.400 ;
    RECT 459.620 1.400 460.460 736.400 ;
    RECT 460.740 1.400 461.580 736.400 ;
    RECT 461.860 1.400 462.700 736.400 ;
    RECT 462.980 1.400 463.820 736.400 ;
    RECT 464.100 1.400 464.940 736.400 ;
    RECT 465.220 1.400 466.060 736.400 ;
    RECT 466.340 1.400 467.180 736.400 ;
    RECT 467.460 1.400 468.300 736.400 ;
    RECT 468.580 1.400 469.420 736.400 ;
    RECT 469.700 1.400 470.540 736.400 ;
    RECT 470.820 1.400 471.660 736.400 ;
    RECT 471.940 1.400 472.780 736.400 ;
    RECT 473.060 1.400 473.900 736.400 ;
    RECT 474.180 1.400 475.020 736.400 ;
    RECT 475.300 1.400 476.140 736.400 ;
    RECT 476.420 1.400 477.260 736.400 ;
    RECT 477.540 1.400 478.380 736.400 ;
    RECT 478.660 1.400 479.500 736.400 ;
    RECT 479.780 1.400 480.620 736.400 ;
    RECT 480.900 1.400 481.740 736.400 ;
    RECT 482.020 1.400 482.860 736.400 ;
    RECT 483.140 1.400 483.980 736.400 ;
    RECT 484.260 1.400 485.100 736.400 ;
    RECT 485.380 1.400 486.220 736.400 ;
    RECT 486.500 1.400 487.340 736.400 ;
    RECT 487.620 1.400 488.460 736.400 ;
    RECT 488.740 1.400 489.580 736.400 ;
    RECT 489.860 1.400 490.700 736.400 ;
    RECT 490.980 1.400 491.820 736.400 ;
    RECT 492.100 1.400 492.940 736.400 ;
    RECT 493.220 1.400 494.060 736.400 ;
    RECT 494.340 1.400 495.180 736.400 ;
    RECT 495.460 1.400 496.300 736.400 ;
    RECT 496.580 1.400 497.420 736.400 ;
    RECT 497.700 1.400 498.540 736.400 ;
    RECT 498.820 1.400 499.660 736.400 ;
    RECT 499.940 1.400 500.780 736.400 ;
    RECT 501.060 1.400 501.900 736.400 ;
    RECT 502.180 1.400 503.020 736.400 ;
    RECT 503.300 1.400 504.140 736.400 ;
    RECT 504.420 1.400 505.260 736.400 ;
    RECT 505.540 1.400 506.380 736.400 ;
    RECT 506.660 1.400 507.500 736.400 ;
    RECT 507.780 1.400 508.620 736.400 ;
    RECT 508.900 1.400 509.740 736.400 ;
    RECT 510.020 1.400 510.860 736.400 ;
    RECT 511.140 1.400 511.980 736.400 ;
    RECT 512.260 1.400 513.100 736.400 ;
    RECT 513.380 1.400 514.220 736.400 ;
    RECT 514.500 1.400 515.340 736.400 ;
    RECT 515.620 1.400 516.460 736.400 ;
    RECT 516.740 1.400 517.580 736.400 ;
    RECT 517.860 1.400 518.700 736.400 ;
    RECT 518.980 1.400 519.820 736.400 ;
    RECT 520.100 1.400 520.940 736.400 ;
    RECT 521.220 1.400 522.060 736.400 ;
    RECT 522.340 1.400 523.180 736.400 ;
    RECT 523.460 1.400 524.300 736.400 ;
    RECT 524.580 1.400 525.420 736.400 ;
    RECT 525.700 1.400 526.540 736.400 ;
    RECT 526.820 1.400 527.660 736.400 ;
    RECT 527.940 1.400 528.780 736.400 ;
    RECT 529.060 1.400 529.900 736.400 ;
    RECT 530.180 1.400 531.020 736.400 ;
    RECT 531.300 1.400 532.140 736.400 ;
    RECT 532.420 1.400 533.260 736.400 ;
    RECT 533.540 1.400 534.380 736.400 ;
    RECT 534.660 1.400 535.500 736.400 ;
    RECT 535.780 1.400 536.620 736.400 ;
    RECT 536.900 1.400 537.740 736.400 ;
    RECT 538.020 1.400 538.860 736.400 ;
    RECT 539.140 1.400 539.980 736.400 ;
    RECT 540.260 1.400 541.100 736.400 ;
    RECT 541.380 1.400 542.220 736.400 ;
    RECT 542.500 1.400 543.340 736.400 ;
    RECT 543.620 1.400 544.460 736.400 ;
    RECT 544.740 1.400 545.580 736.400 ;
    RECT 545.860 1.400 546.700 736.400 ;
    RECT 546.980 1.400 547.820 736.400 ;
    RECT 548.100 1.400 548.940 736.400 ;
    RECT 549.220 1.400 550.060 736.400 ;
    RECT 550.340 1.400 551.180 736.400 ;
    RECT 551.460 1.400 552.300 736.400 ;
    RECT 552.580 1.400 553.420 736.400 ;
    RECT 553.700 1.400 554.540 736.400 ;
    RECT 554.820 1.400 555.660 736.400 ;
    RECT 555.940 1.400 556.780 736.400 ;
    RECT 557.060 1.400 557.900 736.400 ;
    RECT 558.180 1.400 559.020 736.400 ;
    RECT 559.300 1.400 560.140 736.400 ;
    RECT 560.420 1.400 561.260 736.400 ;
    RECT 561.540 1.400 562.380 736.400 ;
    RECT 562.660 1.400 563.500 736.400 ;
    RECT 563.780 1.400 564.620 736.400 ;
    RECT 564.900 1.400 565.740 736.400 ;
    RECT 566.020 1.400 566.860 736.400 ;
    RECT 567.140 1.400 567.980 736.400 ;
    RECT 568.260 1.400 569.100 736.400 ;
    RECT 569.380 1.400 570.220 736.400 ;
    RECT 570.500 1.400 571.340 736.400 ;
    RECT 571.620 1.400 572.460 736.400 ;
    RECT 572.740 1.400 573.580 736.400 ;
    RECT 573.860 1.400 574.700 736.400 ;
    RECT 574.980 1.400 575.820 736.400 ;
    RECT 576.100 1.400 576.940 736.400 ;
    RECT 577.220 1.400 578.060 736.400 ;
    RECT 578.340 1.400 579.180 736.400 ;
    RECT 579.460 1.400 580.300 736.400 ;
    RECT 580.580 1.400 581.420 736.400 ;
    RECT 581.700 1.400 582.540 736.400 ;
    RECT 582.820 1.400 583.660 736.400 ;
    RECT 583.940 1.400 584.780 736.400 ;
    RECT 585.060 1.400 585.900 736.400 ;
    RECT 586.180 1.400 587.020 736.400 ;
    RECT 587.300 1.400 588.140 736.400 ;
    RECT 588.420 1.400 589.260 736.400 ;
    RECT 589.540 1.400 590.380 736.400 ;
    RECT 590.660 1.400 591.500 736.400 ;
    RECT 591.780 1.400 592.620 736.400 ;
    RECT 592.900 1.400 593.740 736.400 ;
    RECT 594.020 1.400 594.860 736.400 ;
    RECT 595.140 1.400 595.980 736.400 ;
    RECT 596.260 1.400 597.100 736.400 ;
    RECT 597.380 1.400 598.220 736.400 ;
    RECT 598.500 1.400 599.340 736.400 ;
    RECT 599.620 1.400 600.460 736.400 ;
    RECT 600.740 1.400 601.580 736.400 ;
    RECT 601.860 1.400 602.700 736.400 ;
    RECT 602.980 1.400 603.820 736.400 ;
    RECT 604.100 1.400 604.940 736.400 ;
    RECT 605.220 1.400 606.060 736.400 ;
    RECT 606.340 1.400 607.180 736.400 ;
    RECT 607.460 1.400 608.300 736.400 ;
    RECT 608.580 1.400 609.420 736.400 ;
    RECT 609.700 1.400 610.540 736.400 ;
    RECT 610.820 1.400 611.660 736.400 ;
    RECT 611.940 1.400 612.780 736.400 ;
    RECT 613.060 1.400 613.900 736.400 ;
    RECT 614.180 1.400 615.020 736.400 ;
    RECT 615.300 1.400 616.140 736.400 ;
    RECT 616.420 1.400 617.260 736.400 ;
    RECT 617.540 1.400 618.380 736.400 ;
    RECT 618.660 1.400 619.500 736.400 ;
    RECT 619.780 1.400 620.620 736.400 ;
    RECT 620.900 1.400 621.740 736.400 ;
    RECT 622.020 1.400 622.860 736.400 ;
    RECT 623.140 1.400 623.980 736.400 ;
    RECT 624.260 1.400 625.100 736.400 ;
    RECT 625.380 1.400 626.220 736.400 ;
    RECT 626.500 1.400 627.340 736.400 ;
    RECT 627.620 1.400 628.460 736.400 ;
    RECT 628.740 1.400 629.580 736.400 ;
    RECT 629.860 1.400 630.700 736.400 ;
    RECT 630.980 1.400 631.820 736.400 ;
    RECT 632.100 1.400 632.940 736.400 ;
    RECT 633.220 1.400 634.060 736.400 ;
    RECT 634.340 1.400 635.180 736.400 ;
    RECT 635.460 1.400 636.300 736.400 ;
    RECT 636.580 1.400 637.420 736.400 ;
    RECT 637.700 1.400 638.540 736.400 ;
    RECT 638.820 1.400 639.660 736.400 ;
    RECT 639.940 1.400 640.780 736.400 ;
    RECT 641.060 1.400 641.900 736.400 ;
    RECT 642.180 1.400 643.020 736.400 ;
    RECT 643.300 1.400 644.140 736.400 ;
    RECT 644.420 1.400 645.260 736.400 ;
    RECT 645.540 1.400 646.380 736.400 ;
    RECT 646.660 1.400 647.500 736.400 ;
    RECT 647.780 1.400 648.620 736.400 ;
    RECT 648.900 1.400 649.740 736.400 ;
    RECT 650.020 1.400 650.860 736.400 ;
    RECT 651.140 1.400 651.980 736.400 ;
    RECT 652.260 1.400 653.100 736.400 ;
    RECT 653.380 1.400 654.220 736.400 ;
    RECT 654.500 1.400 655.340 736.400 ;
    RECT 655.620 1.400 656.460 736.400 ;
    RECT 656.740 1.400 657.580 736.400 ;
    RECT 657.860 1.400 658.700 736.400 ;
    RECT 658.980 1.400 659.820 736.400 ;
    RECT 660.100 1.400 660.940 736.400 ;
    RECT 661.220 1.400 662.060 736.400 ;
    RECT 662.340 1.400 663.180 736.400 ;
    RECT 663.460 1.400 664.300 736.400 ;
    RECT 664.580 1.400 665.420 736.400 ;
    RECT 665.700 1.400 666.540 736.400 ;
    RECT 666.820 1.400 667.660 736.400 ;
    RECT 667.940 1.400 668.780 736.400 ;
    RECT 669.060 1.400 669.900 736.400 ;
    RECT 670.180 1.400 671.020 736.400 ;
    RECT 671.300 1.400 672.140 736.400 ;
    RECT 672.420 1.400 673.260 736.400 ;
    RECT 673.540 1.400 674.380 736.400 ;
    RECT 674.660 1.400 675.500 736.400 ;
    RECT 675.780 1.400 676.620 736.400 ;
    RECT 676.900 1.400 677.740 736.400 ;
    RECT 678.020 1.400 678.860 736.400 ;
    RECT 679.140 1.400 679.980 736.400 ;
    RECT 680.260 1.400 681.100 736.400 ;
    RECT 681.380 1.400 682.220 736.400 ;
    RECT 682.500 1.400 683.340 736.400 ;
    RECT 683.620 1.400 684.460 736.400 ;
    RECT 684.740 1.400 685.580 736.400 ;
    RECT 685.860 1.400 686.700 736.400 ;
    RECT 686.980 1.400 687.820 736.400 ;
    RECT 688.100 1.400 688.940 736.400 ;
    RECT 689.220 1.400 690.060 736.400 ;
    RECT 690.340 1.400 691.180 736.400 ;
    RECT 691.460 1.400 692.300 736.400 ;
    RECT 692.580 1.400 693.420 736.400 ;
    RECT 693.700 1.400 694.540 736.400 ;
    RECT 694.820 1.400 695.660 736.400 ;
    RECT 695.940 1.400 696.780 736.400 ;
    RECT 697.060 1.400 697.900 736.400 ;
    RECT 698.180 1.400 699.020 736.400 ;
    RECT 699.300 1.400 700.140 736.400 ;
    RECT 700.420 1.400 701.260 736.400 ;
    RECT 701.540 1.400 702.380 736.400 ;
    RECT 702.660 1.400 703.500 736.400 ;
    RECT 703.780 1.400 704.620 736.400 ;
    RECT 704.900 1.400 705.740 736.400 ;
    RECT 706.020 1.400 706.860 736.400 ;
    RECT 707.140 1.400 707.980 736.400 ;
    RECT 708.260 1.400 709.100 736.400 ;
    RECT 709.380 1.400 710.220 736.400 ;
    RECT 710.500 1.400 711.340 736.400 ;
    RECT 711.620 1.400 712.460 736.400 ;
    RECT 712.740 1.400 713.580 736.400 ;
    RECT 713.860 1.400 714.700 736.400 ;
    RECT 714.980 1.400 715.820 736.400 ;
    RECT 716.100 1.400 716.940 736.400 ;
    RECT 717.220 1.400 718.060 736.400 ;
    RECT 718.340 1.400 719.180 736.400 ;
    RECT 719.460 1.400 720.300 736.400 ;
    RECT 720.580 1.400 721.420 736.400 ;
    RECT 721.700 1.400 722.540 736.400 ;
    RECT 722.820 1.400 723.660 736.400 ;
    RECT 723.940 1.400 724.780 736.400 ;
    RECT 725.060 1.400 725.900 736.400 ;
    RECT 726.180 1.400 727.020 736.400 ;
    RECT 727.300 1.400 728.140 736.400 ;
    RECT 728.420 1.400 729.260 736.400 ;
    RECT 729.540 1.400 730.380 736.400 ;
    RECT 730.660 1.400 731.500 736.400 ;
    RECT 731.780 1.400 732.620 736.400 ;
    RECT 732.900 1.400 733.740 736.400 ;
    RECT 734.020 1.400 734.860 736.400 ;
    RECT 735.140 1.400 735.980 736.400 ;
    RECT 736.260 1.400 737.100 736.400 ;
    RECT 737.380 1.400 738.220 736.400 ;
    RECT 738.500 1.400 739.340 736.400 ;
    RECT 739.620 1.400 740.460 736.400 ;
    RECT 740.740 1.400 741.580 736.400 ;
    RECT 741.860 1.400 742.700 736.400 ;
    RECT 742.980 1.400 743.820 736.400 ;
    RECT 744.100 1.400 744.940 736.400 ;
    RECT 745.220 1.400 746.060 736.400 ;
    RECT 746.340 1.400 747.180 736.400 ;
    RECT 747.460 1.400 748.300 736.400 ;
    RECT 748.580 1.400 749.420 736.400 ;
    RECT 749.700 1.400 750.540 736.400 ;
    RECT 750.820 1.400 751.660 736.400 ;
    RECT 751.940 1.400 752.780 736.400 ;
    RECT 753.060 1.400 753.900 736.400 ;
    RECT 754.180 1.400 755.020 736.400 ;
    RECT 755.300 1.400 756.140 736.400 ;
    RECT 756.420 1.400 757.260 736.400 ;
    RECT 757.540 1.400 758.380 736.400 ;
    RECT 758.660 1.400 759.500 736.400 ;
    RECT 759.780 1.400 760.620 736.400 ;
    RECT 760.900 1.400 761.740 736.400 ;
    RECT 762.020 1.400 762.860 736.400 ;
    RECT 763.140 1.400 763.980 736.400 ;
    RECT 764.260 1.400 765.100 736.400 ;
    RECT 765.380 1.400 766.220 736.400 ;
    RECT 766.500 1.400 767.340 736.400 ;
    RECT 767.620 1.400 768.460 736.400 ;
    RECT 768.740 1.400 769.580 736.400 ;
    RECT 769.860 1.400 770.700 736.400 ;
    RECT 770.980 1.400 771.820 736.400 ;
    RECT 772.100 1.400 772.940 736.400 ;
    RECT 773.220 1.400 774.060 736.400 ;
    RECT 774.340 1.400 775.180 736.400 ;
    RECT 775.460 1.400 776.300 736.400 ;
    RECT 776.580 1.400 777.420 736.400 ;
    RECT 777.700 1.400 778.540 736.400 ;
    RECT 778.820 1.400 779.660 736.400 ;
    RECT 779.940 1.400 780.780 736.400 ;
    RECT 781.060 1.400 781.900 736.400 ;
    RECT 782.180 1.400 783.020 736.400 ;
    RECT 783.300 1.400 784.140 736.400 ;
    RECT 784.420 1.400 785.260 736.400 ;
    RECT 785.540 1.400 786.380 736.400 ;
    RECT 786.660 1.400 787.500 736.400 ;
    RECT 787.780 1.400 788.620 736.400 ;
    RECT 788.900 1.400 789.740 736.400 ;
    RECT 790.020 1.400 790.860 736.400 ;
    RECT 791.140 1.400 791.980 736.400 ;
    RECT 792.260 1.400 793.100 736.400 ;
    RECT 793.380 1.400 794.220 736.400 ;
    RECT 794.500 1.400 795.340 736.400 ;
    RECT 795.620 1.400 796.460 736.400 ;
    RECT 796.740 1.400 797.580 736.400 ;
    RECT 797.860 1.400 798.700 736.400 ;
    RECT 798.980 1.400 799.820 736.400 ;
    RECT 800.100 1.400 800.940 736.400 ;
    RECT 801.220 1.400 802.060 736.400 ;
    RECT 802.340 1.400 803.180 736.400 ;
    RECT 803.460 1.400 804.300 736.400 ;
    RECT 804.580 1.400 805.420 736.400 ;
    RECT 805.700 1.400 806.540 736.400 ;
    RECT 806.820 1.400 807.660 736.400 ;
    RECT 807.940 1.400 808.780 736.400 ;
    RECT 809.060 1.400 809.900 736.400 ;
    RECT 810.180 1.400 811.020 736.400 ;
    RECT 811.300 1.400 812.140 736.400 ;
    RECT 812.420 1.400 813.260 736.400 ;
    RECT 813.540 1.400 814.380 736.400 ;
    RECT 814.660 1.400 815.500 736.400 ;
    RECT 815.780 1.400 816.620 736.400 ;
    RECT 816.900 1.400 817.740 736.400 ;
    RECT 818.020 1.400 818.860 736.400 ;
    RECT 819.140 1.400 819.980 736.400 ;
    RECT 820.260 1.400 821.100 736.400 ;
    RECT 821.380 1.400 822.220 736.400 ;
    RECT 822.500 1.400 823.340 736.400 ;
    RECT 823.620 1.400 824.460 736.400 ;
    RECT 824.740 1.400 825.580 736.400 ;
    RECT 825.860 1.400 826.700 736.400 ;
    RECT 826.980 1.400 827.820 736.400 ;
    RECT 828.100 1.400 828.940 736.400 ;
    RECT 829.220 1.400 830.060 736.400 ;
    RECT 830.340 1.400 831.180 736.400 ;
    RECT 831.460 1.400 832.300 736.400 ;
    RECT 832.580 1.400 833.420 736.400 ;
    RECT 833.700 1.400 834.540 736.400 ;
    RECT 834.820 1.400 835.660 736.400 ;
    RECT 835.940 1.400 836.780 736.400 ;
    RECT 837.060 1.400 837.900 736.400 ;
    RECT 838.180 1.400 839.020 736.400 ;
    RECT 839.300 1.400 840.140 736.400 ;
    RECT 840.420 1.400 841.260 736.400 ;
    RECT 841.540 1.400 842.380 736.400 ;
    RECT 842.660 1.400 843.500 736.400 ;
    RECT 843.780 1.400 844.620 736.400 ;
    RECT 844.900 1.400 845.740 736.400 ;
    RECT 846.020 1.400 846.860 736.400 ;
    RECT 847.140 1.400 847.980 736.400 ;
    RECT 848.260 1.400 849.100 736.400 ;
    RECT 849.380 1.400 850.220 736.400 ;
    RECT 850.500 1.400 851.340 736.400 ;
    RECT 851.620 1.400 852.460 736.400 ;
    RECT 852.740 1.400 853.580 736.400 ;
    RECT 853.860 1.400 854.700 736.400 ;
    RECT 854.980 1.400 855.820 736.400 ;
    RECT 856.100 1.400 856.940 736.400 ;
    RECT 857.220 1.400 858.060 736.400 ;
    RECT 858.340 1.400 859.180 736.400 ;
    RECT 859.460 1.400 860.300 736.400 ;
    RECT 860.580 1.400 861.420 736.400 ;
    RECT 861.700 1.400 862.540 736.400 ;
    RECT 862.820 1.400 863.660 736.400 ;
    RECT 863.940 1.400 864.780 736.400 ;
    RECT 865.060 1.400 865.900 736.400 ;
    RECT 866.180 1.400 867.020 736.400 ;
    RECT 867.300 1.400 868.140 736.400 ;
    RECT 868.420 1.400 869.260 736.400 ;
    RECT 869.540 1.400 870.380 736.400 ;
    RECT 870.660 1.400 871.500 736.400 ;
    RECT 871.780 1.400 872.620 736.400 ;
    RECT 872.900 1.400 873.740 736.400 ;
    RECT 874.020 1.400 874.860 736.400 ;
    RECT 875.140 1.400 875.980 736.400 ;
    RECT 876.260 1.400 877.100 736.400 ;
    RECT 877.380 1.400 878.220 736.400 ;
    RECT 878.500 1.400 879.340 736.400 ;
    RECT 879.620 1.400 880.460 736.400 ;
    RECT 880.740 1.400 881.580 736.400 ;
    RECT 881.860 1.400 882.700 736.400 ;
    RECT 882.980 1.400 883.820 736.400 ;
    RECT 884.100 1.400 884.940 736.400 ;
    RECT 885.220 1.400 886.060 736.400 ;
    RECT 886.340 1.400 887.180 736.400 ;
    RECT 887.460 1.400 888.300 736.400 ;
    RECT 888.580 1.400 889.420 736.400 ;
    RECT 889.700 1.400 890.540 736.400 ;
    RECT 890.820 1.400 891.660 736.400 ;
    RECT 891.940 1.400 892.780 736.400 ;
    RECT 893.060 1.400 893.900 736.400 ;
    RECT 894.180 1.400 895.020 736.400 ;
    RECT 895.300 1.400 896.140 736.400 ;
    RECT 896.420 1.400 897.260 736.400 ;
    RECT 897.540 1.400 898.380 736.400 ;
    RECT 898.660 1.400 899.500 736.400 ;
    RECT 899.780 1.400 900.620 736.400 ;
    RECT 900.900 1.400 901.740 736.400 ;
    RECT 902.020 1.400 902.860 736.400 ;
    RECT 903.140 1.400 903.980 736.400 ;
    RECT 904.260 1.400 905.100 736.400 ;
    RECT 905.380 1.400 906.220 736.400 ;
    RECT 906.500 1.400 907.340 736.400 ;
    RECT 907.620 1.400 908.460 736.400 ;
    RECT 908.740 1.400 909.580 736.400 ;
    RECT 909.860 1.400 910.700 736.400 ;
    RECT 910.980 1.400 911.820 736.400 ;
    RECT 912.100 1.400 912.940 736.400 ;
    RECT 913.220 1.400 914.060 736.400 ;
    RECT 914.340 1.400 915.180 736.400 ;
    RECT 915.460 1.400 916.300 736.400 ;
    RECT 916.580 1.400 917.420 736.400 ;
    RECT 917.700 1.400 918.540 736.400 ;
    RECT 918.820 1.400 919.660 736.400 ;
    RECT 919.940 1.400 920.780 736.400 ;
    RECT 921.060 1.400 921.900 736.400 ;
    RECT 922.180 1.400 923.020 736.400 ;
    RECT 923.300 1.400 924.140 736.400 ;
    RECT 924.420 1.400 925.260 736.400 ;
    RECT 925.540 1.400 926.380 736.400 ;
    RECT 926.660 1.400 927.500 736.400 ;
    RECT 927.780 1.400 928.620 736.400 ;
    RECT 928.900 1.400 929.740 736.400 ;
    RECT 930.020 1.400 930.860 736.400 ;
    RECT 931.140 1.400 931.980 736.400 ;
    RECT 932.260 1.400 933.100 736.400 ;
    RECT 933.380 1.400 934.220 736.400 ;
    RECT 934.500 1.400 935.340 736.400 ;
    RECT 935.620 1.400 936.460 736.400 ;
    RECT 936.740 1.400 937.580 736.400 ;
    RECT 937.860 1.400 938.700 736.400 ;
    RECT 938.980 1.400 939.820 736.400 ;
    RECT 940.100 1.400 940.940 736.400 ;
    RECT 941.220 1.400 942.060 736.400 ;
    RECT 942.340 1.400 943.180 736.400 ;
    RECT 943.460 1.400 944.300 736.400 ;
    RECT 944.580 1.400 945.420 736.400 ;
    RECT 945.700 1.400 946.540 736.400 ;
    RECT 946.820 1.400 947.660 736.400 ;
    RECT 947.940 1.400 948.780 736.400 ;
    RECT 949.060 1.400 949.900 736.400 ;
    RECT 950.180 1.400 951.020 736.400 ;
    RECT 951.300 1.400 952.140 736.400 ;
    RECT 952.420 1.400 953.260 736.400 ;
    RECT 953.540 1.400 954.380 736.400 ;
    RECT 954.660 1.400 955.500 736.400 ;
    RECT 955.780 1.400 956.620 736.400 ;
    RECT 956.900 1.400 957.740 736.400 ;
    RECT 958.020 1.400 958.860 736.400 ;
    RECT 959.140 1.400 959.980 736.400 ;
    RECT 960.260 1.400 961.100 736.400 ;
    RECT 961.380 1.400 962.220 736.400 ;
    RECT 962.500 1.400 963.340 736.400 ;
    RECT 963.620 1.400 964.460 736.400 ;
    RECT 964.740 1.400 965.580 736.400 ;
    RECT 965.860 1.400 966.700 736.400 ;
    RECT 966.980 1.400 967.820 736.400 ;
    RECT 968.100 1.400 968.940 736.400 ;
    RECT 969.220 1.400 970.060 736.400 ;
    RECT 970.340 1.400 971.180 736.400 ;
    RECT 971.460 1.400 972.300 736.400 ;
    RECT 972.580 1.400 973.420 736.400 ;
    RECT 973.700 1.400 974.540 736.400 ;
    RECT 974.820 1.400 975.660 736.400 ;
    RECT 975.940 1.400 976.780 736.400 ;
    RECT 977.060 1.400 977.900 736.400 ;
    RECT 978.180 1.400 979.020 736.400 ;
    RECT 979.300 1.400 980.140 736.400 ;
    RECT 980.420 1.400 981.260 736.400 ;
    RECT 981.540 1.400 982.380 736.400 ;
    RECT 982.660 1.400 983.500 736.400 ;
    RECT 983.780 1.400 984.620 736.400 ;
    RECT 984.900 1.400 985.740 736.400 ;
    RECT 986.020 1.400 986.860 736.400 ;
    RECT 987.140 1.400 987.980 736.400 ;
    RECT 988.260 1.400 989.100 736.400 ;
    RECT 989.380 1.400 990.220 736.400 ;
    RECT 990.500 1.400 991.340 736.400 ;
    RECT 991.620 1.400 992.460 736.400 ;
    RECT 992.740 1.400 993.580 736.400 ;
    RECT 993.860 1.400 994.700 736.400 ;
    RECT 994.980 1.400 995.820 736.400 ;
    RECT 996.100 1.400 996.940 736.400 ;
    RECT 997.220 1.400 998.060 736.400 ;
    RECT 998.340 1.400 999.180 736.400 ;
    RECT 999.460 1.400 1000.300 736.400 ;
    RECT 1000.580 1.400 1001.420 736.400 ;
    RECT 1001.700 1.400 1002.540 736.400 ;
    RECT 1002.820 1.400 1003.660 736.400 ;
    RECT 1003.940 1.400 1004.780 736.400 ;
    RECT 1005.060 1.400 1005.900 736.400 ;
    RECT 1006.180 1.400 1007.020 736.400 ;
    RECT 1007.300 1.400 1008.140 736.400 ;
    RECT 1008.420 1.400 1009.260 736.400 ;
    RECT 1009.540 1.400 1010.380 736.400 ;
    RECT 1010.660 1.400 1011.500 736.400 ;
    RECT 1011.780 1.400 1012.620 736.400 ;
    RECT 1012.900 1.400 1013.740 736.400 ;
    RECT 1014.020 1.400 1014.860 736.400 ;
    RECT 1015.140 1.400 1015.980 736.400 ;
    RECT 1016.260 1.400 1017.100 736.400 ;
    RECT 1017.380 1.400 1018.220 736.400 ;
    RECT 1018.500 1.400 1019.340 736.400 ;
    RECT 1019.620 1.400 1020.460 736.400 ;
    RECT 1020.740 1.400 1021.580 736.400 ;
    RECT 1021.860 1.400 1022.700 736.400 ;
    RECT 1022.980 1.400 1023.820 736.400 ;
    RECT 1024.100 1.400 1024.940 736.400 ;
    RECT 1025.220 1.400 1026.060 736.400 ;
    RECT 1026.340 1.400 1027.180 736.400 ;
    RECT 1027.460 1.400 1028.300 736.400 ;
    RECT 1028.580 1.400 1029.420 736.400 ;
    RECT 1029.700 1.400 1030.540 736.400 ;
    RECT 1030.820 1.400 1031.660 736.400 ;
    RECT 1031.940 1.400 1032.780 736.400 ;
    RECT 1033.060 1.400 1033.900 736.400 ;
    RECT 1034.180 1.400 1035.020 736.400 ;
    RECT 1035.300 1.400 1036.140 736.400 ;
    RECT 1036.420 1.400 1037.260 736.400 ;
    RECT 1037.540 1.400 1038.380 736.400 ;
    RECT 1038.660 1.400 1039.500 736.400 ;
    RECT 1039.780 1.400 1040.620 736.400 ;
    RECT 1040.900 1.400 1041.740 736.400 ;
    RECT 1042.020 1.400 1042.860 736.400 ;
    RECT 1043.140 1.400 1043.980 736.400 ;
    RECT 1044.260 1.400 1045.100 736.400 ;
    RECT 1045.380 1.400 1046.220 736.400 ;
    RECT 1046.500 1.400 1047.340 736.400 ;
    RECT 1047.620 1.400 1048.460 736.400 ;
    RECT 1048.740 1.400 1049.580 736.400 ;
    RECT 1049.860 1.400 1050.700 736.400 ;
    RECT 1050.980 1.400 1051.820 736.400 ;
    RECT 1052.100 1.400 1052.940 736.400 ;
    RECT 1053.220 1.400 1054.060 736.400 ;
    RECT 1054.340 1.400 1055.180 736.400 ;
    RECT 1055.460 1.400 1056.300 736.400 ;
    RECT 1056.580 1.400 1057.420 736.400 ;
    RECT 1057.700 1.400 1058.540 736.400 ;
    RECT 1058.820 1.400 1059.660 736.400 ;
    RECT 1059.940 1.400 1060.780 736.400 ;
    RECT 1061.060 1.400 1061.900 736.400 ;
    RECT 1062.180 1.400 1063.020 736.400 ;
    RECT 1063.300 1.400 1064.140 736.400 ;
    RECT 1064.420 1.400 1065.260 736.400 ;
    RECT 1065.540 1.400 1066.380 736.400 ;
    RECT 1066.660 1.400 1067.500 736.400 ;
    RECT 1067.780 1.400 1068.620 736.400 ;
    RECT 1068.900 1.400 1069.740 736.400 ;
    RECT 1070.020 1.400 1070.860 736.400 ;
    RECT 1071.140 1.400 1071.980 736.400 ;
    RECT 1072.260 1.400 1073.100 736.400 ;
    RECT 1073.380 1.400 1074.220 736.400 ;
    RECT 1074.500 1.400 1075.340 736.400 ;
    RECT 1075.620 1.400 1076.460 736.400 ;
    RECT 1076.740 1.400 1077.580 736.400 ;
    RECT 1077.860 1.400 1078.700 736.400 ;
    RECT 1078.980 1.400 1079.820 736.400 ;
    RECT 1080.100 1.400 1080.940 736.400 ;
    RECT 1081.220 1.400 1082.060 736.400 ;
    RECT 1082.340 1.400 1083.180 736.400 ;
    RECT 1083.460 1.400 1084.300 736.400 ;
    RECT 1084.580 1.400 1085.420 736.400 ;
    RECT 1085.700 1.400 1086.540 736.400 ;
    RECT 1086.820 1.400 1087.660 736.400 ;
    RECT 1087.940 1.400 1088.780 736.400 ;
    RECT 1089.060 1.400 1089.900 736.400 ;
    RECT 1090.180 1.400 1091.020 736.400 ;
    RECT 1091.300 1.400 1092.140 736.400 ;
    RECT 1092.420 1.400 1093.260 736.400 ;
    RECT 1093.540 1.400 1094.380 736.400 ;
    RECT 1094.660 1.400 1095.500 736.400 ;
    RECT 1095.780 1.400 1096.620 736.400 ;
    RECT 1096.900 1.400 1097.740 736.400 ;
    RECT 1098.020 1.400 1098.860 736.400 ;
    RECT 1099.140 1.400 1099.980 736.400 ;
    RECT 1100.260 1.400 1101.100 736.400 ;
    RECT 1101.380 1.400 1102.220 736.400 ;
    RECT 1102.500 1.400 1103.340 736.400 ;
    RECT 1103.620 1.400 1104.460 736.400 ;
    RECT 1104.740 1.400 1105.580 736.400 ;
    RECT 1105.860 1.400 1106.700 736.400 ;
    RECT 1106.980 1.400 1107.820 736.400 ;
    RECT 1108.100 1.400 1108.940 736.400 ;
    RECT 1109.220 1.400 1110.060 736.400 ;
    RECT 1110.340 1.400 1111.180 736.400 ;
    RECT 1111.460 1.400 1112.300 736.400 ;
    RECT 1112.580 1.400 1113.420 736.400 ;
    RECT 1113.700 1.400 1114.540 736.400 ;
    RECT 1114.820 1.400 1115.660 736.400 ;
    RECT 1115.940 1.400 1116.780 736.400 ;
    RECT 1117.060 1.400 1117.900 736.400 ;
    RECT 1118.180 1.400 1119.020 736.400 ;
    RECT 1119.300 1.400 1120.140 736.400 ;
    RECT 1120.420 1.400 1121.260 736.400 ;
    RECT 1121.540 1.400 1122.380 736.400 ;
    RECT 1122.660 1.400 1123.500 736.400 ;
    RECT 1123.780 1.400 1124.620 736.400 ;
    RECT 1124.900 1.400 1125.740 736.400 ;
    RECT 1126.020 1.400 1126.860 736.400 ;
    RECT 1127.140 1.400 1127.980 736.400 ;
    RECT 1128.260 1.400 1129.100 736.400 ;
    RECT 1129.380 1.400 1130.220 736.400 ;
    RECT 1130.500 1.400 1131.340 736.400 ;
    RECT 1131.620 1.400 1132.460 736.400 ;
    RECT 1132.740 1.400 1133.580 736.400 ;
    RECT 1133.860 1.400 1134.700 736.400 ;
    RECT 1134.980 1.400 1135.820 736.400 ;
    RECT 1136.100 1.400 1136.940 736.400 ;
    RECT 1137.220 1.400 1138.060 736.400 ;
    RECT 1138.340 1.400 1139.180 736.400 ;
    RECT 1139.460 1.400 1140.300 736.400 ;
    RECT 1140.580 1.400 1141.420 736.400 ;
    RECT 1141.700 1.400 1142.540 736.400 ;
    RECT 1142.820 1.400 1143.660 736.400 ;
    RECT 1143.940 1.400 1144.780 736.400 ;
    RECT 1145.060 1.400 1145.900 736.400 ;
    RECT 1146.180 1.400 1147.020 736.400 ;
    RECT 1147.300 1.400 1148.140 736.400 ;
    RECT 1148.420 1.400 1149.260 736.400 ;
    RECT 1149.540 1.400 1150.380 736.400 ;
    RECT 1150.660 1.400 1151.500 736.400 ;
    RECT 1151.780 1.400 1152.620 736.400 ;
    RECT 1152.900 1.400 1153.740 736.400 ;
    RECT 1154.020 1.400 1154.860 736.400 ;
    RECT 1155.140 1.400 1155.980 736.400 ;
    RECT 1156.260 1.400 1157.100 736.400 ;
    RECT 1157.380 1.400 1158.220 736.400 ;
    RECT 1158.500 1.400 1159.340 736.400 ;
    RECT 1159.620 1.400 1160.460 736.400 ;
    RECT 1160.740 1.400 1161.580 736.400 ;
    RECT 1161.860 1.400 1162.700 736.400 ;
    RECT 1162.980 1.400 1163.820 736.400 ;
    RECT 1164.100 1.400 1164.940 736.400 ;
    RECT 1165.220 1.400 1166.060 736.400 ;
    RECT 1166.340 1.400 1167.180 736.400 ;
    RECT 1167.460 1.400 1168.300 736.400 ;
    RECT 1168.580 1.400 1169.420 736.400 ;
    RECT 1169.700 1.400 1170.540 736.400 ;
    RECT 1170.820 1.400 1171.660 736.400 ;
    RECT 1171.940 1.400 1172.780 736.400 ;
    RECT 1173.060 1.400 1173.900 736.400 ;
    RECT 1174.180 1.400 1175.020 736.400 ;
    RECT 1175.300 1.400 1176.140 736.400 ;
    RECT 1176.420 1.400 1177.260 736.400 ;
    RECT 1177.540 1.400 1178.380 736.400 ;
    RECT 1178.660 1.400 1179.500 736.400 ;
    RECT 1179.780 1.400 1180.620 736.400 ;
    RECT 1180.900 1.400 1181.740 736.400 ;
    RECT 1182.020 1.400 1182.860 736.400 ;
    RECT 1183.140 1.400 1183.980 736.400 ;
    RECT 1184.260 1.400 1185.100 736.400 ;
    RECT 1185.380 1.400 1186.220 736.400 ;
    RECT 1186.500 1.400 1187.340 736.400 ;
    RECT 1187.620 1.400 1188.460 736.400 ;
    RECT 1188.740 1.400 1189.580 736.400 ;
    RECT 1189.860 1.400 1190.700 736.400 ;
    RECT 1190.980 1.400 1191.820 736.400 ;
    RECT 1192.100 1.400 1192.940 736.400 ;
    RECT 1193.220 1.400 1194.060 736.400 ;
    RECT 1194.340 1.400 1195.180 736.400 ;
    RECT 1195.460 1.400 1196.300 736.400 ;
    RECT 1196.580 1.400 1197.420 736.400 ;
    RECT 1197.700 1.400 1198.540 736.400 ;
    RECT 1198.820 1.400 1199.660 736.400 ;
    RECT 1199.940 1.400 1200.780 736.400 ;
    RECT 1201.060 1.400 1201.900 736.400 ;
    RECT 1202.180 1.400 1203.020 736.400 ;
    RECT 1203.300 1.400 1204.140 736.400 ;
    RECT 1204.420 1.400 1205.260 736.400 ;
    RECT 1205.540 1.400 1206.380 736.400 ;
    RECT 1206.660 1.400 1207.500 736.400 ;
    RECT 1207.780 1.400 1208.620 736.400 ;
    RECT 1208.900 1.400 1209.740 736.400 ;
    RECT 1210.020 1.400 1210.860 736.400 ;
    RECT 1211.140 1.400 1211.980 736.400 ;
    RECT 1212.260 1.400 1213.100 736.400 ;
    RECT 1213.380 1.400 1214.220 736.400 ;
    RECT 1214.500 1.400 1215.340 736.400 ;
    RECT 1215.620 1.400 1216.460 736.400 ;
    RECT 1216.740 1.400 1217.580 736.400 ;
    RECT 1217.860 1.400 1218.700 736.400 ;
    RECT 1218.980 1.400 1219.820 736.400 ;
    RECT 1220.100 1.400 1220.940 736.400 ;
    RECT 1221.220 1.400 1222.060 736.400 ;
    RECT 1222.340 1.400 1223.180 736.400 ;
    RECT 1223.460 1.400 1224.300 736.400 ;
    RECT 1224.580 1.400 1225.420 736.400 ;
    RECT 1225.700 1.400 1226.540 736.400 ;
    RECT 1226.820 1.400 1227.660 736.400 ;
    RECT 1227.940 1.400 1228.780 736.400 ;
    RECT 1229.060 1.400 1229.900 736.400 ;
    RECT 1230.180 1.400 1231.020 736.400 ;
    RECT 1231.300 1.400 1232.140 736.400 ;
    RECT 1232.420 1.400 1233.260 736.400 ;
    RECT 1233.540 1.400 1234.380 736.400 ;
    RECT 1234.660 1.400 1235.500 736.400 ;
    RECT 1235.780 1.400 1236.620 736.400 ;
    RECT 1236.900 1.400 1237.740 736.400 ;
    RECT 1238.020 1.400 1238.860 736.400 ;
    RECT 1239.140 1.400 1239.980 736.400 ;
    RECT 1240.260 1.400 1241.100 736.400 ;
    RECT 1241.380 1.400 1242.220 736.400 ;
    RECT 1242.500 1.400 1243.340 736.400 ;
    RECT 1243.620 1.400 1244.460 736.400 ;
    RECT 1244.740 1.400 1245.580 736.400 ;
    RECT 1245.860 1.400 1246.700 736.400 ;
    RECT 1246.980 1.400 1247.820 736.400 ;
    RECT 1248.100 1.400 1248.940 736.400 ;
    RECT 1249.220 1.400 1250.060 736.400 ;
    RECT 1250.340 1.400 1251.180 736.400 ;
    RECT 1251.460 1.400 1252.300 736.400 ;
    RECT 1252.580 1.400 1253.420 736.400 ;
    RECT 1253.700 1.400 1254.540 736.400 ;
    RECT 1254.820 1.400 1255.660 736.400 ;
    RECT 1255.940 1.400 1256.780 736.400 ;
    RECT 1257.060 1.400 1257.900 736.400 ;
    RECT 1258.180 1.400 1259.020 736.400 ;
    RECT 1259.300 1.400 1260.140 736.400 ;
    RECT 1260.420 1.400 1261.260 736.400 ;
    RECT 1261.540 1.400 1262.380 736.400 ;
    RECT 1262.660 1.400 1263.500 736.400 ;
    RECT 1263.780 1.400 1264.620 736.400 ;
    RECT 1264.900 1.400 1265.740 736.400 ;
    RECT 1266.020 1.400 1266.860 736.400 ;
    RECT 1267.140 1.400 1267.980 736.400 ;
    RECT 1268.260 1.400 1269.100 736.400 ;
    RECT 1269.380 1.400 1270.220 736.400 ;
    RECT 1270.500 1.400 1271.340 736.400 ;
    RECT 1271.620 1.400 1272.460 736.400 ;
    RECT 1272.740 1.400 1273.580 736.400 ;
    RECT 1273.860 1.400 1274.700 736.400 ;
    RECT 1274.980 1.400 1275.820 736.400 ;
    RECT 1276.100 1.400 1276.940 736.400 ;
    RECT 1277.220 1.400 1278.060 736.400 ;
    RECT 1278.340 1.400 1279.180 736.400 ;
    RECT 1279.460 1.400 1280.300 736.400 ;
    RECT 1280.580 1.400 1281.420 736.400 ;
    RECT 1281.700 1.400 1282.540 736.400 ;
    RECT 1282.820 1.400 1283.660 736.400 ;
    RECT 1283.940 1.400 1284.780 736.400 ;
    RECT 1285.060 1.400 1285.900 736.400 ;
    RECT 1286.180 1.400 1287.020 736.400 ;
    RECT 1287.300 1.400 1288.140 736.400 ;
    RECT 1288.420 1.400 1289.260 736.400 ;
    RECT 1289.540 1.400 1290.380 736.400 ;
    RECT 1290.660 1.400 1291.500 736.400 ;
    RECT 1291.780 1.400 1292.620 736.400 ;
    RECT 1292.900 1.400 1293.740 736.400 ;
    RECT 1294.020 1.400 1294.860 736.400 ;
    RECT 1295.140 1.400 1295.980 736.400 ;
    RECT 1296.260 1.400 1297.100 736.400 ;
    RECT 1297.380 1.400 1298.220 736.400 ;
    RECT 1298.500 1.400 1299.340 736.400 ;
    RECT 1299.620 1.400 1300.460 736.400 ;
    RECT 1300.740 1.400 1301.580 736.400 ;
    RECT 1301.860 1.400 1302.700 736.400 ;
    RECT 1302.980 1.400 1303.820 736.400 ;
    RECT 1304.100 1.400 1304.940 736.400 ;
    RECT 1305.220 1.400 1306.060 736.400 ;
    RECT 1306.340 1.400 1307.180 736.400 ;
    RECT 1307.460 1.400 1308.300 736.400 ;
    RECT 1308.580 1.400 1309.420 736.400 ;
    RECT 1309.700 1.400 1310.540 736.400 ;
    RECT 1310.820 1.400 1311.660 736.400 ;
    RECT 1311.940 1.400 1312.780 736.400 ;
    RECT 1313.060 1.400 1313.900 736.400 ;
    RECT 1314.180 1.400 1315.020 736.400 ;
    RECT 1315.300 1.400 1316.140 736.400 ;
    RECT 1316.420 1.400 1317.260 736.400 ;
    RECT 1317.540 1.400 1318.380 736.400 ;
    RECT 1318.660 1.400 1319.500 736.400 ;
    RECT 1319.780 1.400 1320.620 736.400 ;
    RECT 1320.900 1.400 1321.740 736.400 ;
    RECT 1322.020 1.400 1322.860 736.400 ;
    RECT 1323.140 1.400 1323.980 736.400 ;
    RECT 1324.260 1.400 1325.100 736.400 ;
    RECT 1325.380 1.400 1326.220 736.400 ;
    RECT 1326.500 1.400 1327.340 736.400 ;
    RECT 1327.620 1.400 1328.460 736.400 ;
    RECT 1328.740 1.400 1329.580 736.400 ;
    RECT 1329.860 1.400 1330.700 736.400 ;
    RECT 1330.980 1.400 1331.820 736.400 ;
    RECT 1332.100 1.400 1332.940 736.400 ;
    RECT 1333.220 1.400 1334.060 736.400 ;
    RECT 1334.340 1.400 1335.180 736.400 ;
    RECT 1335.460 1.400 1336.300 736.400 ;
    RECT 1336.580 1.400 1337.420 736.400 ;
    RECT 1337.700 1.400 1338.540 736.400 ;
    RECT 1338.820 1.400 1339.660 736.400 ;
    RECT 1339.940 1.400 1340.780 736.400 ;
    RECT 1341.060 1.400 1341.900 736.400 ;
    RECT 1342.180 1.400 1343.020 736.400 ;
    RECT 1343.300 1.400 1344.140 736.400 ;
    RECT 1344.420 1.400 1345.260 736.400 ;
    RECT 1345.540 1.400 1346.380 736.400 ;
    RECT 1346.660 1.400 1347.500 736.400 ;
    RECT 1347.780 1.400 1348.620 736.400 ;
    RECT 1348.900 1.400 1349.740 736.400 ;
    RECT 1350.020 1.400 1350.860 736.400 ;
    RECT 1351.140 1.400 1351.980 736.400 ;
    RECT 1352.260 1.400 1353.100 736.400 ;
    RECT 1353.380 1.400 1354.220 736.400 ;
    RECT 1354.500 1.400 1355.340 736.400 ;
    RECT 1355.620 1.400 1356.460 736.400 ;
    RECT 1356.740 1.400 1357.580 736.400 ;
    RECT 1357.860 1.400 1358.700 736.400 ;
    RECT 1358.980 1.400 1359.820 736.400 ;
    RECT 1360.100 1.400 1360.940 736.400 ;
    RECT 1361.220 1.400 1362.060 736.400 ;
    RECT 1362.340 1.400 1363.180 736.400 ;
    RECT 1363.460 1.400 1364.300 736.400 ;
    RECT 1364.580 1.400 1365.420 736.400 ;
    RECT 1365.700 1.400 1366.540 736.400 ;
    RECT 1366.820 1.400 1367.660 736.400 ;
    RECT 1367.940 1.400 1368.780 736.400 ;
    RECT 1369.060 1.400 1369.900 736.400 ;
    RECT 1370.180 1.400 1371.020 736.400 ;
    RECT 1371.300 1.400 1372.140 736.400 ;
    RECT 1372.420 1.400 1373.260 736.400 ;
    RECT 1373.540 1.400 1374.380 736.400 ;
    RECT 1374.660 1.400 1375.500 736.400 ;
    RECT 1375.780 1.400 1376.620 736.400 ;
    RECT 1376.900 1.400 1377.740 736.400 ;
    RECT 1378.020 1.400 1378.860 736.400 ;
    RECT 1379.140 1.400 1379.980 736.400 ;
    RECT 1380.260 1.400 1381.100 736.400 ;
    RECT 1381.380 1.400 1382.220 736.400 ;
    RECT 1382.500 1.400 1383.340 736.400 ;
    RECT 1383.620 1.400 1384.460 736.400 ;
    RECT 1384.740 1.400 1385.580 736.400 ;
    RECT 1385.860 1.400 1386.700 736.400 ;
    RECT 1386.980 1.400 1387.820 736.400 ;
    RECT 1388.100 1.400 1388.940 736.400 ;
    RECT 1389.220 1.400 1390.060 736.400 ;
    RECT 1390.340 1.400 1391.180 736.400 ;
    RECT 1391.460 1.400 1392.300 736.400 ;
    RECT 1392.580 1.400 1393.420 736.400 ;
    RECT 1393.700 1.400 1394.540 736.400 ;
    RECT 1394.820 1.400 1395.660 736.400 ;
    RECT 1395.940 1.400 1396.780 736.400 ;
    RECT 1397.060 1.400 1397.900 736.400 ;
    RECT 1398.180 1.400 1399.020 736.400 ;
    RECT 1399.300 1.400 1400.140 736.400 ;
    RECT 1400.420 1.400 1401.260 736.400 ;
    RECT 1401.540 1.400 1402.380 736.400 ;
    RECT 1402.660 1.400 1403.500 736.400 ;
    RECT 1403.780 1.400 1404.620 736.400 ;
    RECT 1404.900 1.400 1405.740 736.400 ;
    RECT 1406.020 1.400 1406.860 736.400 ;
    RECT 1407.140 1.400 1407.980 736.400 ;
    RECT 1408.260 1.400 1409.100 736.400 ;
    RECT 1409.380 1.400 1410.220 736.400 ;
    RECT 1410.500 1.400 1411.340 736.400 ;
    RECT 1411.620 1.400 1412.460 736.400 ;
    RECT 1412.740 1.400 1413.580 736.400 ;
    RECT 1413.860 1.400 1414.700 736.400 ;
    RECT 1414.980 1.400 1415.820 736.400 ;
    RECT 1416.100 1.400 1416.940 736.400 ;
    RECT 1417.220 1.400 1418.060 736.400 ;
    RECT 1418.340 1.400 1419.180 736.400 ;
    RECT 1419.460 1.400 1420.300 736.400 ;
    RECT 1420.580 1.400 1421.420 736.400 ;
    RECT 1421.700 1.400 1422.540 736.400 ;
    RECT 1422.820 1.400 1423.660 736.400 ;
    RECT 1423.940 1.400 1424.780 736.400 ;
    RECT 1425.060 1.400 1425.900 736.400 ;
    RECT 1426.180 1.400 1427.020 736.400 ;
    RECT 1427.300 1.400 1428.140 736.400 ;
    RECT 1428.420 1.400 1429.260 736.400 ;
    RECT 1429.540 1.400 1430.380 736.400 ;
    RECT 1430.660 1.400 1431.500 736.400 ;
    RECT 1431.780 1.400 1432.620 736.400 ;
    RECT 1432.900 1.400 1433.740 736.400 ;
    RECT 1434.020 1.400 1434.860 736.400 ;
    RECT 1435.140 1.400 1435.980 736.400 ;
    RECT 1436.260 1.400 1437.100 736.400 ;
    RECT 1437.380 1.400 1438.220 736.400 ;
    RECT 1438.500 1.400 1439.340 736.400 ;
    RECT 1439.620 1.400 1440.460 736.400 ;
    RECT 1440.740 1.400 1441.580 736.400 ;
    RECT 1441.860 1.400 1442.700 736.400 ;
    RECT 1442.980 1.400 1443.820 736.400 ;
    RECT 1444.100 1.400 1444.940 736.400 ;
    RECT 1445.220 1.400 1446.060 736.400 ;
    RECT 1446.340 1.400 1447.180 736.400 ;
    RECT 1447.460 1.400 1448.300 736.400 ;
    RECT 1448.580 1.400 1449.420 736.400 ;
    RECT 1449.700 1.400 1450.540 736.400 ;
    RECT 1450.820 1.400 1451.660 736.400 ;
    RECT 1451.940 1.400 1452.780 736.400 ;
    RECT 1453.060 1.400 1453.900 736.400 ;
    RECT 1454.180 1.400 1455.020 736.400 ;
    RECT 1455.300 1.400 1456.140 736.400 ;
    RECT 1456.420 1.400 1457.260 736.400 ;
    RECT 1457.540 1.400 1458.380 736.400 ;
    RECT 1458.660 1.400 1459.500 736.400 ;
    RECT 1459.780 1.400 1460.620 736.400 ;
    RECT 1460.900 1.400 1461.740 736.400 ;
    RECT 1462.020 1.400 1462.860 736.400 ;
    RECT 1463.140 1.400 1463.980 736.400 ;
    RECT 1464.260 1.400 1465.100 736.400 ;
    RECT 1465.380 1.400 1466.220 736.400 ;
    RECT 1466.500 1.400 1467.340 736.400 ;
    RECT 1467.620 1.400 1468.460 736.400 ;
    RECT 1468.740 1.400 1469.580 736.400 ;
    RECT 1469.860 1.400 1470.700 736.400 ;
    RECT 1470.980 1.400 1471.820 736.400 ;
    RECT 1472.100 1.400 1472.940 736.400 ;
    RECT 1473.220 1.400 1474.060 736.400 ;
    RECT 1474.340 1.400 1475.180 736.400 ;
    RECT 1475.460 1.400 1476.300 736.400 ;
    RECT 1476.580 1.400 1477.420 736.400 ;
    RECT 1477.700 1.400 1478.540 736.400 ;
    RECT 1478.820 1.400 1479.660 736.400 ;
    RECT 1479.940 1.400 1480.780 736.400 ;
    RECT 1481.060 1.400 1481.900 736.400 ;
    RECT 1482.180 1.400 1483.020 736.400 ;
    RECT 1483.300 1.400 1484.140 736.400 ;
    RECT 1484.420 1.400 1485.260 736.400 ;
    RECT 1485.540 1.400 1486.380 736.400 ;
    RECT 1486.660 1.400 1487.500 736.400 ;
    RECT 1487.780 1.400 1488.620 736.400 ;
    RECT 1488.900 1.400 1489.740 736.400 ;
    RECT 1490.020 1.400 1490.860 736.400 ;
    RECT 1491.140 1.400 1491.980 736.400 ;
    RECT 1492.260 1.400 1493.100 736.400 ;
    RECT 1493.380 1.400 1494.220 736.400 ;
    RECT 1494.500 1.400 1495.340 736.400 ;
    RECT 1495.620 1.400 1496.460 736.400 ;
    RECT 1496.740 1.400 1497.580 736.400 ;
    RECT 1497.860 1.400 1498.700 736.400 ;
    RECT 1498.980 1.400 1499.820 736.400 ;
    RECT 1500.100 1.400 1500.940 736.400 ;
    RECT 1501.220 1.400 1502.060 736.400 ;
    RECT 1502.340 1.400 1503.180 736.400 ;
    RECT 1503.460 1.400 1504.300 736.400 ;
    RECT 1504.580 1.400 1505.420 736.400 ;
    RECT 1505.700 1.400 1506.540 736.400 ;
    RECT 1506.820 1.400 1507.660 736.400 ;
    RECT 1507.940 1.400 1508.780 736.400 ;
    RECT 1509.060 1.400 1509.900 736.400 ;
    RECT 1510.180 1.400 1511.020 736.400 ;
    RECT 1511.300 1.400 1512.140 736.400 ;
    RECT 1512.420 1.400 1513.260 736.400 ;
    RECT 1513.540 1.400 1514.380 736.400 ;
    RECT 1514.660 1.400 1515.500 736.400 ;
    RECT 1515.780 1.400 1516.620 736.400 ;
    RECT 1516.900 1.400 1517.740 736.400 ;
    RECT 1518.020 1.400 1518.860 736.400 ;
    RECT 1519.140 1.400 1519.980 736.400 ;
    RECT 1520.260 1.400 1521.100 736.400 ;
    RECT 1521.380 1.400 1522.220 736.400 ;
    RECT 1522.500 1.400 1523.340 736.400 ;
    RECT 1523.620 1.400 1524.460 736.400 ;
    RECT 1524.740 1.400 1525.580 736.400 ;
    RECT 1525.860 1.400 1526.700 736.400 ;
    RECT 1526.980 1.400 1527.820 736.400 ;
    RECT 1528.100 1.400 1528.940 736.400 ;
    RECT 1529.220 1.400 1530.060 736.400 ;
    RECT 1530.340 1.400 1531.180 736.400 ;
    RECT 1531.460 1.400 1532.300 736.400 ;
    RECT 1532.580 1.400 1533.420 736.400 ;
    RECT 1533.700 1.400 1534.540 736.400 ;
    RECT 1534.820 1.400 1535.660 736.400 ;
    RECT 1535.940 1.400 1536.780 736.400 ;
    RECT 1537.060 1.400 1537.900 736.400 ;
    RECT 1538.180 1.400 1539.020 736.400 ;
    RECT 1539.300 1.400 1540.140 736.400 ;
    RECT 1540.420 1.400 1541.260 736.400 ;
    RECT 1541.540 1.400 1542.380 736.400 ;
    RECT 1542.660 1.400 1543.500 736.400 ;
    RECT 1543.780 1.400 1544.620 736.400 ;
    RECT 1544.900 1.400 1545.740 736.400 ;
    RECT 1546.020 1.400 1546.860 736.400 ;
    RECT 1547.140 1.400 1547.980 736.400 ;
    RECT 1548.260 1.400 1549.100 736.400 ;
    RECT 1549.380 1.400 1550.220 736.400 ;
    RECT 1550.500 1.400 1551.340 736.400 ;
    RECT 1551.620 1.400 1552.460 736.400 ;
    RECT 1552.740 1.400 1553.580 736.400 ;
    RECT 1553.860 1.400 1554.700 736.400 ;
    RECT 1554.980 1.400 1555.820 736.400 ;
    RECT 1556.100 1.400 1556.940 736.400 ;
    RECT 1557.220 1.400 1558.060 736.400 ;
    RECT 1558.340 1.400 1559.180 736.400 ;
    RECT 1559.460 1.400 1560.300 736.400 ;
    RECT 1560.580 1.400 1561.420 736.400 ;
    RECT 1561.700 1.400 1562.540 736.400 ;
    RECT 1562.820 1.400 1563.660 736.400 ;
    RECT 1563.940 1.400 1564.780 736.400 ;
    RECT 1565.060 1.400 1565.900 736.400 ;
    RECT 1566.180 1.400 1567.020 736.400 ;
    RECT 1567.300 1.400 1568.140 736.400 ;
    RECT 1568.420 1.400 1569.260 736.400 ;
    RECT 1569.540 1.400 1570.380 736.400 ;
    RECT 1570.660 1.400 1571.500 736.400 ;
    RECT 1571.780 1.400 1572.620 736.400 ;
    RECT 1572.900 1.400 1573.740 736.400 ;
    RECT 1574.020 1.400 1574.860 736.400 ;
    RECT 1575.140 1.400 1575.980 736.400 ;
    RECT 1576.260 1.400 1577.100 736.400 ;
    RECT 1577.380 1.400 1578.220 736.400 ;
    RECT 1578.500 1.400 1579.340 736.400 ;
    RECT 1579.620 1.400 1580.460 736.400 ;
    RECT 1580.740 1.400 1581.580 736.400 ;
    RECT 1581.860 1.400 1582.700 736.400 ;
    RECT 1582.980 1.400 1583.820 736.400 ;
    RECT 1584.100 1.400 1584.940 736.400 ;
    RECT 1585.220 1.400 1586.060 736.400 ;
    RECT 1586.340 1.400 1587.180 736.400 ;
    RECT 1587.460 1.400 1588.300 736.400 ;
    RECT 1588.580 1.400 1589.420 736.400 ;
    RECT 1589.700 1.400 1590.540 736.400 ;
    RECT 1590.820 1.400 1591.660 736.400 ;
    RECT 1591.940 1.400 1592.780 736.400 ;
    RECT 1593.060 1.400 1593.900 736.400 ;
    RECT 1594.180 1.400 1595.020 736.400 ;
    RECT 1595.300 1.400 1596.140 736.400 ;
    RECT 1596.420 1.400 1597.260 736.400 ;
    RECT 1597.540 1.400 1598.380 736.400 ;
    RECT 1598.660 1.400 1599.500 736.400 ;
    RECT 1599.780 1.400 1600.620 736.400 ;
    RECT 1600.900 1.400 1601.740 736.400 ;
    RECT 1602.020 1.400 1602.860 736.400 ;
    RECT 1603.140 1.400 1603.980 736.400 ;
    RECT 1604.260 1.400 1605.100 736.400 ;
    RECT 1605.380 1.400 1606.220 736.400 ;
    RECT 1606.500 1.400 1607.340 736.400 ;
    RECT 1607.620 1.400 1608.460 736.400 ;
    RECT 1608.740 1.400 1609.580 736.400 ;
    RECT 1609.860 1.400 1610.700 736.400 ;
    RECT 1610.980 1.400 1611.820 736.400 ;
    RECT 1612.100 1.400 1612.940 736.400 ;
    RECT 1613.220 1.400 1614.060 736.400 ;
    RECT 1614.340 1.400 1615.180 736.400 ;
    RECT 1615.460 1.400 1616.300 736.400 ;
    RECT 1616.580 1.400 1617.420 736.400 ;
    RECT 1617.700 1.400 1618.540 736.400 ;
    RECT 1618.820 1.400 1619.660 736.400 ;
    RECT 1619.940 1.400 1620.780 736.400 ;
    RECT 1621.060 1.400 1621.900 736.400 ;
    RECT 1622.180 1.400 1623.020 736.400 ;
    RECT 1623.300 1.400 1624.140 736.400 ;
    RECT 1624.420 1.400 1625.260 736.400 ;
    RECT 1625.540 1.400 1626.380 736.400 ;
    RECT 1626.660 1.400 1627.500 736.400 ;
    RECT 1627.780 1.400 1628.620 736.400 ;
    RECT 1628.900 1.400 1629.740 736.400 ;
    RECT 1630.020 1.400 1631.530 736.400 ;
    LAYER OVERLAP ;
    RECT 0 0 1631.530 737.800 ;
  END
END sram_256x4096_1rw

END LIBRARY
