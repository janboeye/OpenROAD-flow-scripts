VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_512x4096_1rw
  FOREIGN sram_512x4096_1rw 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 2064.540 BY 1281.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.865 0.070 4.935 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.065 0.070 9.135 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.265 0.070 13.335 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.465 0.070 17.535 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.665 0.070 21.735 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.665 0.070 28.735 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.065 0.070 30.135 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.865 0.070 32.935 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.265 0.070 34.335 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.365 0.070 36.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.465 0.070 38.535 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.665 0.070 42.735 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.665 0.070 49.735 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.065 0.070 51.135 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.165 0.070 53.235 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.865 0.070 53.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.265 0.070 55.335 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.065 0.070 58.135 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.465 0.070 59.535 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.565 0.070 61.635 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.265 0.070 62.335 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.665 0.070 63.735 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.465 0.070 66.535 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.865 0.070 67.935 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.665 0.070 70.735 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.065 0.070 72.135 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.865 0.070 74.935 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.265 0.070 76.335 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.065 0.070 79.135 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.465 0.070 80.535 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.265 0.070 83.335 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.665 0.070 84.735 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.465 0.070 87.535 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.865 0.070 88.935 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.965 0.070 91.035 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.665 0.070 91.735 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.065 0.070 93.135 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.765 0.070 93.835 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.165 0.070 95.235 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.865 0.070 95.935 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.265 0.070 97.335 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.965 0.070 98.035 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.665 0.070 98.735 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.365 0.070 99.435 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.065 0.070 100.135 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.465 0.070 101.535 ;
    END
  END w_mask_in[143]
  PIN w_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.165 0.070 102.235 ;
    END
  END w_mask_in[144]
  PIN w_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.865 0.070 102.935 ;
    END
  END w_mask_in[145]
  PIN w_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.565 0.070 103.635 ;
    END
  END w_mask_in[146]
  PIN w_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.265 0.070 104.335 ;
    END
  END w_mask_in[147]
  PIN w_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.965 0.070 105.035 ;
    END
  END w_mask_in[148]
  PIN w_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.665 0.070 105.735 ;
    END
  END w_mask_in[149]
  PIN w_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.365 0.070 106.435 ;
    END
  END w_mask_in[150]
  PIN w_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.065 0.070 107.135 ;
    END
  END w_mask_in[151]
  PIN w_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.765 0.070 107.835 ;
    END
  END w_mask_in[152]
  PIN w_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.465 0.070 108.535 ;
    END
  END w_mask_in[153]
  PIN w_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END w_mask_in[154]
  PIN w_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.865 0.070 109.935 ;
    END
  END w_mask_in[155]
  PIN w_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.565 0.070 110.635 ;
    END
  END w_mask_in[156]
  PIN w_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.265 0.070 111.335 ;
    END
  END w_mask_in[157]
  PIN w_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.965 0.070 112.035 ;
    END
  END w_mask_in[158]
  PIN w_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.665 0.070 112.735 ;
    END
  END w_mask_in[159]
  PIN w_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.365 0.070 113.435 ;
    END
  END w_mask_in[160]
  PIN w_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.065 0.070 114.135 ;
    END
  END w_mask_in[161]
  PIN w_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.765 0.070 114.835 ;
    END
  END w_mask_in[162]
  PIN w_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.465 0.070 115.535 ;
    END
  END w_mask_in[163]
  PIN w_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END w_mask_in[164]
  PIN w_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.865 0.070 116.935 ;
    END
  END w_mask_in[165]
  PIN w_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END w_mask_in[166]
  PIN w_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.265 0.070 118.335 ;
    END
  END w_mask_in[167]
  PIN w_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END w_mask_in[168]
  PIN w_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.665 0.070 119.735 ;
    END
  END w_mask_in[169]
  PIN w_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.365 0.070 120.435 ;
    END
  END w_mask_in[170]
  PIN w_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.065 0.070 121.135 ;
    END
  END w_mask_in[171]
  PIN w_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.765 0.070 121.835 ;
    END
  END w_mask_in[172]
  PIN w_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.465 0.070 122.535 ;
    END
  END w_mask_in[173]
  PIN w_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.165 0.070 123.235 ;
    END
  END w_mask_in[174]
  PIN w_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.865 0.070 123.935 ;
    END
  END w_mask_in[175]
  PIN w_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.565 0.070 124.635 ;
    END
  END w_mask_in[176]
  PIN w_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.265 0.070 125.335 ;
    END
  END w_mask_in[177]
  PIN w_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.965 0.070 126.035 ;
    END
  END w_mask_in[178]
  PIN w_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.665 0.070 126.735 ;
    END
  END w_mask_in[179]
  PIN w_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.365 0.070 127.435 ;
    END
  END w_mask_in[180]
  PIN w_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.065 0.070 128.135 ;
    END
  END w_mask_in[181]
  PIN w_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END w_mask_in[182]
  PIN w_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.465 0.070 129.535 ;
    END
  END w_mask_in[183]
  PIN w_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.165 0.070 130.235 ;
    END
  END w_mask_in[184]
  PIN w_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.865 0.070 130.935 ;
    END
  END w_mask_in[185]
  PIN w_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.565 0.070 131.635 ;
    END
  END w_mask_in[186]
  PIN w_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.265 0.070 132.335 ;
    END
  END w_mask_in[187]
  PIN w_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.965 0.070 133.035 ;
    END
  END w_mask_in[188]
  PIN w_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.665 0.070 133.735 ;
    END
  END w_mask_in[189]
  PIN w_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.365 0.070 134.435 ;
    END
  END w_mask_in[190]
  PIN w_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.065 0.070 135.135 ;
    END
  END w_mask_in[191]
  PIN w_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.765 0.070 135.835 ;
    END
  END w_mask_in[192]
  PIN w_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.465 0.070 136.535 ;
    END
  END w_mask_in[193]
  PIN w_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.165 0.070 137.235 ;
    END
  END w_mask_in[194]
  PIN w_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.865 0.070 137.935 ;
    END
  END w_mask_in[195]
  PIN w_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.565 0.070 138.635 ;
    END
  END w_mask_in[196]
  PIN w_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.265 0.070 139.335 ;
    END
  END w_mask_in[197]
  PIN w_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END w_mask_in[198]
  PIN w_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.665 0.070 140.735 ;
    END
  END w_mask_in[199]
  PIN w_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.365 0.070 141.435 ;
    END
  END w_mask_in[200]
  PIN w_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.065 0.070 142.135 ;
    END
  END w_mask_in[201]
  PIN w_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.765 0.070 142.835 ;
    END
  END w_mask_in[202]
  PIN w_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.465 0.070 143.535 ;
    END
  END w_mask_in[203]
  PIN w_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.165 0.070 144.235 ;
    END
  END w_mask_in[204]
  PIN w_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.865 0.070 144.935 ;
    END
  END w_mask_in[205]
  PIN w_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.565 0.070 145.635 ;
    END
  END w_mask_in[206]
  PIN w_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.265 0.070 146.335 ;
    END
  END w_mask_in[207]
  PIN w_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.965 0.070 147.035 ;
    END
  END w_mask_in[208]
  PIN w_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.665 0.070 147.735 ;
    END
  END w_mask_in[209]
  PIN w_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END w_mask_in[210]
  PIN w_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.065 0.070 149.135 ;
    END
  END w_mask_in[211]
  PIN w_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.765 0.070 149.835 ;
    END
  END w_mask_in[212]
  PIN w_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.465 0.070 150.535 ;
    END
  END w_mask_in[213]
  PIN w_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.165 0.070 151.235 ;
    END
  END w_mask_in[214]
  PIN w_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.865 0.070 151.935 ;
    END
  END w_mask_in[215]
  PIN w_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.565 0.070 152.635 ;
    END
  END w_mask_in[216]
  PIN w_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.265 0.070 153.335 ;
    END
  END w_mask_in[217]
  PIN w_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.965 0.070 154.035 ;
    END
  END w_mask_in[218]
  PIN w_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.665 0.070 154.735 ;
    END
  END w_mask_in[219]
  PIN w_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.365 0.070 155.435 ;
    END
  END w_mask_in[220]
  PIN w_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.065 0.070 156.135 ;
    END
  END w_mask_in[221]
  PIN w_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.765 0.070 156.835 ;
    END
  END w_mask_in[222]
  PIN w_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.465 0.070 157.535 ;
    END
  END w_mask_in[223]
  PIN w_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.165 0.070 158.235 ;
    END
  END w_mask_in[224]
  PIN w_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.865 0.070 158.935 ;
    END
  END w_mask_in[225]
  PIN w_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.565 0.070 159.635 ;
    END
  END w_mask_in[226]
  PIN w_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.265 0.070 160.335 ;
    END
  END w_mask_in[227]
  PIN w_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.965 0.070 161.035 ;
    END
  END w_mask_in[228]
  PIN w_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.665 0.070 161.735 ;
    END
  END w_mask_in[229]
  PIN w_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.365 0.070 162.435 ;
    END
  END w_mask_in[230]
  PIN w_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.065 0.070 163.135 ;
    END
  END w_mask_in[231]
  PIN w_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.765 0.070 163.835 ;
    END
  END w_mask_in[232]
  PIN w_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.465 0.070 164.535 ;
    END
  END w_mask_in[233]
  PIN w_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END w_mask_in[234]
  PIN w_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.865 0.070 165.935 ;
    END
  END w_mask_in[235]
  PIN w_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.565 0.070 166.635 ;
    END
  END w_mask_in[236]
  PIN w_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.265 0.070 167.335 ;
    END
  END w_mask_in[237]
  PIN w_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.965 0.070 168.035 ;
    END
  END w_mask_in[238]
  PIN w_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.665 0.070 168.735 ;
    END
  END w_mask_in[239]
  PIN w_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.365 0.070 169.435 ;
    END
  END w_mask_in[240]
  PIN w_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.065 0.070 170.135 ;
    END
  END w_mask_in[241]
  PIN w_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.765 0.070 170.835 ;
    END
  END w_mask_in[242]
  PIN w_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.465 0.070 171.535 ;
    END
  END w_mask_in[243]
  PIN w_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END w_mask_in[244]
  PIN w_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.865 0.070 172.935 ;
    END
  END w_mask_in[245]
  PIN w_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.565 0.070 173.635 ;
    END
  END w_mask_in[246]
  PIN w_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.265 0.070 174.335 ;
    END
  END w_mask_in[247]
  PIN w_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.965 0.070 175.035 ;
    END
  END w_mask_in[248]
  PIN w_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.665 0.070 175.735 ;
    END
  END w_mask_in[249]
  PIN w_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.365 0.070 176.435 ;
    END
  END w_mask_in[250]
  PIN w_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.065 0.070 177.135 ;
    END
  END w_mask_in[251]
  PIN w_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END w_mask_in[252]
  PIN w_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.465 0.070 178.535 ;
    END
  END w_mask_in[253]
  PIN w_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.165 0.070 179.235 ;
    END
  END w_mask_in[254]
  PIN w_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.865 0.070 179.935 ;
    END
  END w_mask_in[255]
  PIN w_mask_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.565 0.070 180.635 ;
    END
  END w_mask_in[256]
  PIN w_mask_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.265 0.070 181.335 ;
    END
  END w_mask_in[257]
  PIN w_mask_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.965 0.070 182.035 ;
    END
  END w_mask_in[258]
  PIN w_mask_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.665 0.070 182.735 ;
    END
  END w_mask_in[259]
  PIN w_mask_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.365 0.070 183.435 ;
    END
  END w_mask_in[260]
  PIN w_mask_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.065 0.070 184.135 ;
    END
  END w_mask_in[261]
  PIN w_mask_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.765 0.070 184.835 ;
    END
  END w_mask_in[262]
  PIN w_mask_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.465 0.070 185.535 ;
    END
  END w_mask_in[263]
  PIN w_mask_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.165 0.070 186.235 ;
    END
  END w_mask_in[264]
  PIN w_mask_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.865 0.070 186.935 ;
    END
  END w_mask_in[265]
  PIN w_mask_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.565 0.070 187.635 ;
    END
  END w_mask_in[266]
  PIN w_mask_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.265 0.070 188.335 ;
    END
  END w_mask_in[267]
  PIN w_mask_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.965 0.070 189.035 ;
    END
  END w_mask_in[268]
  PIN w_mask_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.665 0.070 189.735 ;
    END
  END w_mask_in[269]
  PIN w_mask_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.365 0.070 190.435 ;
    END
  END w_mask_in[270]
  PIN w_mask_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.065 0.070 191.135 ;
    END
  END w_mask_in[271]
  PIN w_mask_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.765 0.070 191.835 ;
    END
  END w_mask_in[272]
  PIN w_mask_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.465 0.070 192.535 ;
    END
  END w_mask_in[273]
  PIN w_mask_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.165 0.070 193.235 ;
    END
  END w_mask_in[274]
  PIN w_mask_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.865 0.070 193.935 ;
    END
  END w_mask_in[275]
  PIN w_mask_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.565 0.070 194.635 ;
    END
  END w_mask_in[276]
  PIN w_mask_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.265 0.070 195.335 ;
    END
  END w_mask_in[277]
  PIN w_mask_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.965 0.070 196.035 ;
    END
  END w_mask_in[278]
  PIN w_mask_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.665 0.070 196.735 ;
    END
  END w_mask_in[279]
  PIN w_mask_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END w_mask_in[280]
  PIN w_mask_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.065 0.070 198.135 ;
    END
  END w_mask_in[281]
  PIN w_mask_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.765 0.070 198.835 ;
    END
  END w_mask_in[282]
  PIN w_mask_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.465 0.070 199.535 ;
    END
  END w_mask_in[283]
  PIN w_mask_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.165 0.070 200.235 ;
    END
  END w_mask_in[284]
  PIN w_mask_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.865 0.070 200.935 ;
    END
  END w_mask_in[285]
  PIN w_mask_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.565 0.070 201.635 ;
    END
  END w_mask_in[286]
  PIN w_mask_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.265 0.070 202.335 ;
    END
  END w_mask_in[287]
  PIN w_mask_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.965 0.070 203.035 ;
    END
  END w_mask_in[288]
  PIN w_mask_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.665 0.070 203.735 ;
    END
  END w_mask_in[289]
  PIN w_mask_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.365 0.070 204.435 ;
    END
  END w_mask_in[290]
  PIN w_mask_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.065 0.070 205.135 ;
    END
  END w_mask_in[291]
  PIN w_mask_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.765 0.070 205.835 ;
    END
  END w_mask_in[292]
  PIN w_mask_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.465 0.070 206.535 ;
    END
  END w_mask_in[293]
  PIN w_mask_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.165 0.070 207.235 ;
    END
  END w_mask_in[294]
  PIN w_mask_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.865 0.070 207.935 ;
    END
  END w_mask_in[295]
  PIN w_mask_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.565 0.070 208.635 ;
    END
  END w_mask_in[296]
  PIN w_mask_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.265 0.070 209.335 ;
    END
  END w_mask_in[297]
  PIN w_mask_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.965 0.070 210.035 ;
    END
  END w_mask_in[298]
  PIN w_mask_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.665 0.070 210.735 ;
    END
  END w_mask_in[299]
  PIN w_mask_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.365 0.070 211.435 ;
    END
  END w_mask_in[300]
  PIN w_mask_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.065 0.070 212.135 ;
    END
  END w_mask_in[301]
  PIN w_mask_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.765 0.070 212.835 ;
    END
  END w_mask_in[302]
  PIN w_mask_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.465 0.070 213.535 ;
    END
  END w_mask_in[303]
  PIN w_mask_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.165 0.070 214.235 ;
    END
  END w_mask_in[304]
  PIN w_mask_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.865 0.070 214.935 ;
    END
  END w_mask_in[305]
  PIN w_mask_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.565 0.070 215.635 ;
    END
  END w_mask_in[306]
  PIN w_mask_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.265 0.070 216.335 ;
    END
  END w_mask_in[307]
  PIN w_mask_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.965 0.070 217.035 ;
    END
  END w_mask_in[308]
  PIN w_mask_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.665 0.070 217.735 ;
    END
  END w_mask_in[309]
  PIN w_mask_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.365 0.070 218.435 ;
    END
  END w_mask_in[310]
  PIN w_mask_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.065 0.070 219.135 ;
    END
  END w_mask_in[311]
  PIN w_mask_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.765 0.070 219.835 ;
    END
  END w_mask_in[312]
  PIN w_mask_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.465 0.070 220.535 ;
    END
  END w_mask_in[313]
  PIN w_mask_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.165 0.070 221.235 ;
    END
  END w_mask_in[314]
  PIN w_mask_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.865 0.070 221.935 ;
    END
  END w_mask_in[315]
  PIN w_mask_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.565 0.070 222.635 ;
    END
  END w_mask_in[316]
  PIN w_mask_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.265 0.070 223.335 ;
    END
  END w_mask_in[317]
  PIN w_mask_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.965 0.070 224.035 ;
    END
  END w_mask_in[318]
  PIN w_mask_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.665 0.070 224.735 ;
    END
  END w_mask_in[319]
  PIN w_mask_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.365 0.070 225.435 ;
    END
  END w_mask_in[320]
  PIN w_mask_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.065 0.070 226.135 ;
    END
  END w_mask_in[321]
  PIN w_mask_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END w_mask_in[322]
  PIN w_mask_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.465 0.070 227.535 ;
    END
  END w_mask_in[323]
  PIN w_mask_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.165 0.070 228.235 ;
    END
  END w_mask_in[324]
  PIN w_mask_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.865 0.070 228.935 ;
    END
  END w_mask_in[325]
  PIN w_mask_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.565 0.070 229.635 ;
    END
  END w_mask_in[326]
  PIN w_mask_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.265 0.070 230.335 ;
    END
  END w_mask_in[327]
  PIN w_mask_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.965 0.070 231.035 ;
    END
  END w_mask_in[328]
  PIN w_mask_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.665 0.070 231.735 ;
    END
  END w_mask_in[329]
  PIN w_mask_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.365 0.070 232.435 ;
    END
  END w_mask_in[330]
  PIN w_mask_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.065 0.070 233.135 ;
    END
  END w_mask_in[331]
  PIN w_mask_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.765 0.070 233.835 ;
    END
  END w_mask_in[332]
  PIN w_mask_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.465 0.070 234.535 ;
    END
  END w_mask_in[333]
  PIN w_mask_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.165 0.070 235.235 ;
    END
  END w_mask_in[334]
  PIN w_mask_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.865 0.070 235.935 ;
    END
  END w_mask_in[335]
  PIN w_mask_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.565 0.070 236.635 ;
    END
  END w_mask_in[336]
  PIN w_mask_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.265 0.070 237.335 ;
    END
  END w_mask_in[337]
  PIN w_mask_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.965 0.070 238.035 ;
    END
  END w_mask_in[338]
  PIN w_mask_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.665 0.070 238.735 ;
    END
  END w_mask_in[339]
  PIN w_mask_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.365 0.070 239.435 ;
    END
  END w_mask_in[340]
  PIN w_mask_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.065 0.070 240.135 ;
    END
  END w_mask_in[341]
  PIN w_mask_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.765 0.070 240.835 ;
    END
  END w_mask_in[342]
  PIN w_mask_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.465 0.070 241.535 ;
    END
  END w_mask_in[343]
  PIN w_mask_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.165 0.070 242.235 ;
    END
  END w_mask_in[344]
  PIN w_mask_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.865 0.070 242.935 ;
    END
  END w_mask_in[345]
  PIN w_mask_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.565 0.070 243.635 ;
    END
  END w_mask_in[346]
  PIN w_mask_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.265 0.070 244.335 ;
    END
  END w_mask_in[347]
  PIN w_mask_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.965 0.070 245.035 ;
    END
  END w_mask_in[348]
  PIN w_mask_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.665 0.070 245.735 ;
    END
  END w_mask_in[349]
  PIN w_mask_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.365 0.070 246.435 ;
    END
  END w_mask_in[350]
  PIN w_mask_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.065 0.070 247.135 ;
    END
  END w_mask_in[351]
  PIN w_mask_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.765 0.070 247.835 ;
    END
  END w_mask_in[352]
  PIN w_mask_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.465 0.070 248.535 ;
    END
  END w_mask_in[353]
  PIN w_mask_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.165 0.070 249.235 ;
    END
  END w_mask_in[354]
  PIN w_mask_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.865 0.070 249.935 ;
    END
  END w_mask_in[355]
  PIN w_mask_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.565 0.070 250.635 ;
    END
  END w_mask_in[356]
  PIN w_mask_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.265 0.070 251.335 ;
    END
  END w_mask_in[357]
  PIN w_mask_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.965 0.070 252.035 ;
    END
  END w_mask_in[358]
  PIN w_mask_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.665 0.070 252.735 ;
    END
  END w_mask_in[359]
  PIN w_mask_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.365 0.070 253.435 ;
    END
  END w_mask_in[360]
  PIN w_mask_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.065 0.070 254.135 ;
    END
  END w_mask_in[361]
  PIN w_mask_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.765 0.070 254.835 ;
    END
  END w_mask_in[362]
  PIN w_mask_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.465 0.070 255.535 ;
    END
  END w_mask_in[363]
  PIN w_mask_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.165 0.070 256.235 ;
    END
  END w_mask_in[364]
  PIN w_mask_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.865 0.070 256.935 ;
    END
  END w_mask_in[365]
  PIN w_mask_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.565 0.070 257.635 ;
    END
  END w_mask_in[366]
  PIN w_mask_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.265 0.070 258.335 ;
    END
  END w_mask_in[367]
  PIN w_mask_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.965 0.070 259.035 ;
    END
  END w_mask_in[368]
  PIN w_mask_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.665 0.070 259.735 ;
    END
  END w_mask_in[369]
  PIN w_mask_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.365 0.070 260.435 ;
    END
  END w_mask_in[370]
  PIN w_mask_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.065 0.070 261.135 ;
    END
  END w_mask_in[371]
  PIN w_mask_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.765 0.070 261.835 ;
    END
  END w_mask_in[372]
  PIN w_mask_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.465 0.070 262.535 ;
    END
  END w_mask_in[373]
  PIN w_mask_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.165 0.070 263.235 ;
    END
  END w_mask_in[374]
  PIN w_mask_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.865 0.070 263.935 ;
    END
  END w_mask_in[375]
  PIN w_mask_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.565 0.070 264.635 ;
    END
  END w_mask_in[376]
  PIN w_mask_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.265 0.070 265.335 ;
    END
  END w_mask_in[377]
  PIN w_mask_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.965 0.070 266.035 ;
    END
  END w_mask_in[378]
  PIN w_mask_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.665 0.070 266.735 ;
    END
  END w_mask_in[379]
  PIN w_mask_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.365 0.070 267.435 ;
    END
  END w_mask_in[380]
  PIN w_mask_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.065 0.070 268.135 ;
    END
  END w_mask_in[381]
  PIN w_mask_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.765 0.070 268.835 ;
    END
  END w_mask_in[382]
  PIN w_mask_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.465 0.070 269.535 ;
    END
  END w_mask_in[383]
  PIN w_mask_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.165 0.070 270.235 ;
    END
  END w_mask_in[384]
  PIN w_mask_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.865 0.070 270.935 ;
    END
  END w_mask_in[385]
  PIN w_mask_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.565 0.070 271.635 ;
    END
  END w_mask_in[386]
  PIN w_mask_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.265 0.070 272.335 ;
    END
  END w_mask_in[387]
  PIN w_mask_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.965 0.070 273.035 ;
    END
  END w_mask_in[388]
  PIN w_mask_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.665 0.070 273.735 ;
    END
  END w_mask_in[389]
  PIN w_mask_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.365 0.070 274.435 ;
    END
  END w_mask_in[390]
  PIN w_mask_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.065 0.070 275.135 ;
    END
  END w_mask_in[391]
  PIN w_mask_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.765 0.070 275.835 ;
    END
  END w_mask_in[392]
  PIN w_mask_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.465 0.070 276.535 ;
    END
  END w_mask_in[393]
  PIN w_mask_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.165 0.070 277.235 ;
    END
  END w_mask_in[394]
  PIN w_mask_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.865 0.070 277.935 ;
    END
  END w_mask_in[395]
  PIN w_mask_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.565 0.070 278.635 ;
    END
  END w_mask_in[396]
  PIN w_mask_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.265 0.070 279.335 ;
    END
  END w_mask_in[397]
  PIN w_mask_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.965 0.070 280.035 ;
    END
  END w_mask_in[398]
  PIN w_mask_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.665 0.070 280.735 ;
    END
  END w_mask_in[399]
  PIN w_mask_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.365 0.070 281.435 ;
    END
  END w_mask_in[400]
  PIN w_mask_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.065 0.070 282.135 ;
    END
  END w_mask_in[401]
  PIN w_mask_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.765 0.070 282.835 ;
    END
  END w_mask_in[402]
  PIN w_mask_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.465 0.070 283.535 ;
    END
  END w_mask_in[403]
  PIN w_mask_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.165 0.070 284.235 ;
    END
  END w_mask_in[404]
  PIN w_mask_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.865 0.070 284.935 ;
    END
  END w_mask_in[405]
  PIN w_mask_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.565 0.070 285.635 ;
    END
  END w_mask_in[406]
  PIN w_mask_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.265 0.070 286.335 ;
    END
  END w_mask_in[407]
  PIN w_mask_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.965 0.070 287.035 ;
    END
  END w_mask_in[408]
  PIN w_mask_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.665 0.070 287.735 ;
    END
  END w_mask_in[409]
  PIN w_mask_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.365 0.070 288.435 ;
    END
  END w_mask_in[410]
  PIN w_mask_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.065 0.070 289.135 ;
    END
  END w_mask_in[411]
  PIN w_mask_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.765 0.070 289.835 ;
    END
  END w_mask_in[412]
  PIN w_mask_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.465 0.070 290.535 ;
    END
  END w_mask_in[413]
  PIN w_mask_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.165 0.070 291.235 ;
    END
  END w_mask_in[414]
  PIN w_mask_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.865 0.070 291.935 ;
    END
  END w_mask_in[415]
  PIN w_mask_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.565 0.070 292.635 ;
    END
  END w_mask_in[416]
  PIN w_mask_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.265 0.070 293.335 ;
    END
  END w_mask_in[417]
  PIN w_mask_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.965 0.070 294.035 ;
    END
  END w_mask_in[418]
  PIN w_mask_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.665 0.070 294.735 ;
    END
  END w_mask_in[419]
  PIN w_mask_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.365 0.070 295.435 ;
    END
  END w_mask_in[420]
  PIN w_mask_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.065 0.070 296.135 ;
    END
  END w_mask_in[421]
  PIN w_mask_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.765 0.070 296.835 ;
    END
  END w_mask_in[422]
  PIN w_mask_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.465 0.070 297.535 ;
    END
  END w_mask_in[423]
  PIN w_mask_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.165 0.070 298.235 ;
    END
  END w_mask_in[424]
  PIN w_mask_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.865 0.070 298.935 ;
    END
  END w_mask_in[425]
  PIN w_mask_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.565 0.070 299.635 ;
    END
  END w_mask_in[426]
  PIN w_mask_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.265 0.070 300.335 ;
    END
  END w_mask_in[427]
  PIN w_mask_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.965 0.070 301.035 ;
    END
  END w_mask_in[428]
  PIN w_mask_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.665 0.070 301.735 ;
    END
  END w_mask_in[429]
  PIN w_mask_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.365 0.070 302.435 ;
    END
  END w_mask_in[430]
  PIN w_mask_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.065 0.070 303.135 ;
    END
  END w_mask_in[431]
  PIN w_mask_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.765 0.070 303.835 ;
    END
  END w_mask_in[432]
  PIN w_mask_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.465 0.070 304.535 ;
    END
  END w_mask_in[433]
  PIN w_mask_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.165 0.070 305.235 ;
    END
  END w_mask_in[434]
  PIN w_mask_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.865 0.070 305.935 ;
    END
  END w_mask_in[435]
  PIN w_mask_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.565 0.070 306.635 ;
    END
  END w_mask_in[436]
  PIN w_mask_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.265 0.070 307.335 ;
    END
  END w_mask_in[437]
  PIN w_mask_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.965 0.070 308.035 ;
    END
  END w_mask_in[438]
  PIN w_mask_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.665 0.070 308.735 ;
    END
  END w_mask_in[439]
  PIN w_mask_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.365 0.070 309.435 ;
    END
  END w_mask_in[440]
  PIN w_mask_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.065 0.070 310.135 ;
    END
  END w_mask_in[441]
  PIN w_mask_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.765 0.070 310.835 ;
    END
  END w_mask_in[442]
  PIN w_mask_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.465 0.070 311.535 ;
    END
  END w_mask_in[443]
  PIN w_mask_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.165 0.070 312.235 ;
    END
  END w_mask_in[444]
  PIN w_mask_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.865 0.070 312.935 ;
    END
  END w_mask_in[445]
  PIN w_mask_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.565 0.070 313.635 ;
    END
  END w_mask_in[446]
  PIN w_mask_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.265 0.070 314.335 ;
    END
  END w_mask_in[447]
  PIN w_mask_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.965 0.070 315.035 ;
    END
  END w_mask_in[448]
  PIN w_mask_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.665 0.070 315.735 ;
    END
  END w_mask_in[449]
  PIN w_mask_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.365 0.070 316.435 ;
    END
  END w_mask_in[450]
  PIN w_mask_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.065 0.070 317.135 ;
    END
  END w_mask_in[451]
  PIN w_mask_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.765 0.070 317.835 ;
    END
  END w_mask_in[452]
  PIN w_mask_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.465 0.070 318.535 ;
    END
  END w_mask_in[453]
  PIN w_mask_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.165 0.070 319.235 ;
    END
  END w_mask_in[454]
  PIN w_mask_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.865 0.070 319.935 ;
    END
  END w_mask_in[455]
  PIN w_mask_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.565 0.070 320.635 ;
    END
  END w_mask_in[456]
  PIN w_mask_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.265 0.070 321.335 ;
    END
  END w_mask_in[457]
  PIN w_mask_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.965 0.070 322.035 ;
    END
  END w_mask_in[458]
  PIN w_mask_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.665 0.070 322.735 ;
    END
  END w_mask_in[459]
  PIN w_mask_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.365 0.070 323.435 ;
    END
  END w_mask_in[460]
  PIN w_mask_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.065 0.070 324.135 ;
    END
  END w_mask_in[461]
  PIN w_mask_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.765 0.070 324.835 ;
    END
  END w_mask_in[462]
  PIN w_mask_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.465 0.070 325.535 ;
    END
  END w_mask_in[463]
  PIN w_mask_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.165 0.070 326.235 ;
    END
  END w_mask_in[464]
  PIN w_mask_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.865 0.070 326.935 ;
    END
  END w_mask_in[465]
  PIN w_mask_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.565 0.070 327.635 ;
    END
  END w_mask_in[466]
  PIN w_mask_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.265 0.070 328.335 ;
    END
  END w_mask_in[467]
  PIN w_mask_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.965 0.070 329.035 ;
    END
  END w_mask_in[468]
  PIN w_mask_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.665 0.070 329.735 ;
    END
  END w_mask_in[469]
  PIN w_mask_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.365 0.070 330.435 ;
    END
  END w_mask_in[470]
  PIN w_mask_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.065 0.070 331.135 ;
    END
  END w_mask_in[471]
  PIN w_mask_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.765 0.070 331.835 ;
    END
  END w_mask_in[472]
  PIN w_mask_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.465 0.070 332.535 ;
    END
  END w_mask_in[473]
  PIN w_mask_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.165 0.070 333.235 ;
    END
  END w_mask_in[474]
  PIN w_mask_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.865 0.070 333.935 ;
    END
  END w_mask_in[475]
  PIN w_mask_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.565 0.070 334.635 ;
    END
  END w_mask_in[476]
  PIN w_mask_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.265 0.070 335.335 ;
    END
  END w_mask_in[477]
  PIN w_mask_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.965 0.070 336.035 ;
    END
  END w_mask_in[478]
  PIN w_mask_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.665 0.070 336.735 ;
    END
  END w_mask_in[479]
  PIN w_mask_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.365 0.070 337.435 ;
    END
  END w_mask_in[480]
  PIN w_mask_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.065 0.070 338.135 ;
    END
  END w_mask_in[481]
  PIN w_mask_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.765 0.070 338.835 ;
    END
  END w_mask_in[482]
  PIN w_mask_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.465 0.070 339.535 ;
    END
  END w_mask_in[483]
  PIN w_mask_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.165 0.070 340.235 ;
    END
  END w_mask_in[484]
  PIN w_mask_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.865 0.070 340.935 ;
    END
  END w_mask_in[485]
  PIN w_mask_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.565 0.070 341.635 ;
    END
  END w_mask_in[486]
  PIN w_mask_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.265 0.070 342.335 ;
    END
  END w_mask_in[487]
  PIN w_mask_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.965 0.070 343.035 ;
    END
  END w_mask_in[488]
  PIN w_mask_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.665 0.070 343.735 ;
    END
  END w_mask_in[489]
  PIN w_mask_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.365 0.070 344.435 ;
    END
  END w_mask_in[490]
  PIN w_mask_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.065 0.070 345.135 ;
    END
  END w_mask_in[491]
  PIN w_mask_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.765 0.070 345.835 ;
    END
  END w_mask_in[492]
  PIN w_mask_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.465 0.070 346.535 ;
    END
  END w_mask_in[493]
  PIN w_mask_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.165 0.070 347.235 ;
    END
  END w_mask_in[494]
  PIN w_mask_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.865 0.070 347.935 ;
    END
  END w_mask_in[495]
  PIN w_mask_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.565 0.070 348.635 ;
    END
  END w_mask_in[496]
  PIN w_mask_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.265 0.070 349.335 ;
    END
  END w_mask_in[497]
  PIN w_mask_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.965 0.070 350.035 ;
    END
  END w_mask_in[498]
  PIN w_mask_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.665 0.070 350.735 ;
    END
  END w_mask_in[499]
  PIN w_mask_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.365 0.070 351.435 ;
    END
  END w_mask_in[500]
  PIN w_mask_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.065 0.070 352.135 ;
    END
  END w_mask_in[501]
  PIN w_mask_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.765 0.070 352.835 ;
    END
  END w_mask_in[502]
  PIN w_mask_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.465 0.070 353.535 ;
    END
  END w_mask_in[503]
  PIN w_mask_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.165 0.070 354.235 ;
    END
  END w_mask_in[504]
  PIN w_mask_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.865 0.070 354.935 ;
    END
  END w_mask_in[505]
  PIN w_mask_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.565 0.070 355.635 ;
    END
  END w_mask_in[506]
  PIN w_mask_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.265 0.070 356.335 ;
    END
  END w_mask_in[507]
  PIN w_mask_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.965 0.070 357.035 ;
    END
  END w_mask_in[508]
  PIN w_mask_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.665 0.070 357.735 ;
    END
  END w_mask_in[509]
  PIN w_mask_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.365 0.070 358.435 ;
    END
  END w_mask_in[510]
  PIN w_mask_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.065 0.070 359.135 ;
    END
  END w_mask_in[511]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.085 0.070 407.155 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 407.785 0.070 407.855 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 408.485 0.070 408.555 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 409.185 0.070 409.255 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 409.885 0.070 409.955 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 410.585 0.070 410.655 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.285 0.070 411.355 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.985 0.070 412.055 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 412.685 0.070 412.755 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 413.385 0.070 413.455 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.085 0.070 414.155 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 414.785 0.070 414.855 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 415.485 0.070 415.555 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.185 0.070 416.255 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.885 0.070 416.955 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 417.585 0.070 417.655 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.285 0.070 418.355 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 418.985 0.070 419.055 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.685 0.070 419.755 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 420.385 0.070 420.455 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.085 0.070 421.155 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 421.785 0.070 421.855 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 422.485 0.070 422.555 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.185 0.070 423.255 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 423.885 0.070 423.955 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 424.585 0.070 424.655 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.285 0.070 425.355 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.985 0.070 426.055 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 426.685 0.070 426.755 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.385 0.070 427.455 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.085 0.070 428.155 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.785 0.070 428.855 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 429.485 0.070 429.555 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.185 0.070 430.255 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 430.885 0.070 430.955 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 431.585 0.070 431.655 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.285 0.070 432.355 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.985 0.070 433.055 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 433.685 0.070 433.755 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 434.385 0.070 434.455 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 435.085 0.070 435.155 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 435.785 0.070 435.855 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 436.485 0.070 436.555 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.185 0.070 437.255 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.885 0.070 437.955 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.585 0.070 438.655 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.285 0.070 439.355 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 439.985 0.070 440.055 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 440.685 0.070 440.755 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 441.385 0.070 441.455 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.085 0.070 442.155 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 442.785 0.070 442.855 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.485 0.070 443.555 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.185 0.070 444.255 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 444.885 0.070 444.955 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 445.585 0.070 445.655 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.285 0.070 446.355 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.985 0.070 447.055 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 447.685 0.070 447.755 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.385 0.070 448.455 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.085 0.070 449.155 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.785 0.070 449.855 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 450.485 0.070 450.555 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 451.185 0.070 451.255 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 451.885 0.070 451.955 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 452.585 0.070 452.655 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 453.285 0.070 453.355 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 453.985 0.070 454.055 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.685 0.070 454.755 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 455.385 0.070 455.455 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 456.085 0.070 456.155 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 456.785 0.070 456.855 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 457.485 0.070 457.555 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 458.185 0.070 458.255 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 458.885 0.070 458.955 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 459.585 0.070 459.655 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.285 0.070 460.355 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.985 0.070 461.055 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 461.685 0.070 461.755 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 462.385 0.070 462.455 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 463.085 0.070 463.155 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 463.785 0.070 463.855 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 464.485 0.070 464.555 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.185 0.070 465.255 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 465.885 0.070 465.955 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 466.585 0.070 466.655 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 467.285 0.070 467.355 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 467.985 0.070 468.055 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 468.685 0.070 468.755 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 469.385 0.070 469.455 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.085 0.070 470.155 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.785 0.070 470.855 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 471.485 0.070 471.555 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.185 0.070 472.255 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.885 0.070 472.955 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 473.585 0.070 473.655 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.285 0.070 474.355 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 474.985 0.070 475.055 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.685 0.070 475.755 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 476.385 0.070 476.455 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 477.085 0.070 477.155 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 477.785 0.070 477.855 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 478.485 0.070 478.555 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.185 0.070 479.255 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 479.885 0.070 479.955 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 480.585 0.070 480.655 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.285 0.070 481.355 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.985 0.070 482.055 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 482.685 0.070 482.755 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 483.385 0.070 483.455 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.085 0.070 484.155 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.785 0.070 484.855 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 485.485 0.070 485.555 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.185 0.070 486.255 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.885 0.070 486.955 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 487.585 0.070 487.655 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 488.285 0.070 488.355 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 488.985 0.070 489.055 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 489.685 0.070 489.755 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 490.385 0.070 490.455 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 491.085 0.070 491.155 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 491.785 0.070 491.855 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 492.485 0.070 492.555 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.185 0.070 493.255 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.885 0.070 493.955 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 494.585 0.070 494.655 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 495.285 0.070 495.355 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 495.985 0.070 496.055 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 496.685 0.070 496.755 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 497.385 0.070 497.455 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 498.085 0.070 498.155 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 498.785 0.070 498.855 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 499.485 0.070 499.555 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 500.185 0.070 500.255 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 500.885 0.070 500.955 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 501.585 0.070 501.655 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 502.285 0.070 502.355 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 502.985 0.070 503.055 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 503.685 0.070 503.755 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.385 0.070 504.455 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.085 0.070 505.155 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.785 0.070 505.855 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.485 0.070 506.555 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.185 0.070 507.255 ;
    END
  END rd_out[143]
  PIN rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.885 0.070 507.955 ;
    END
  END rd_out[144]
  PIN rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.585 0.070 508.655 ;
    END
  END rd_out[145]
  PIN rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.285 0.070 509.355 ;
    END
  END rd_out[146]
  PIN rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.985 0.070 510.055 ;
    END
  END rd_out[147]
  PIN rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.685 0.070 510.755 ;
    END
  END rd_out[148]
  PIN rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.385 0.070 511.455 ;
    END
  END rd_out[149]
  PIN rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.085 0.070 512.155 ;
    END
  END rd_out[150]
  PIN rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.785 0.070 512.855 ;
    END
  END rd_out[151]
  PIN rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.485 0.070 513.555 ;
    END
  END rd_out[152]
  PIN rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.185 0.070 514.255 ;
    END
  END rd_out[153]
  PIN rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.885 0.070 514.955 ;
    END
  END rd_out[154]
  PIN rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.585 0.070 515.655 ;
    END
  END rd_out[155]
  PIN rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.285 0.070 516.355 ;
    END
  END rd_out[156]
  PIN rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.985 0.070 517.055 ;
    END
  END rd_out[157]
  PIN rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.685 0.070 517.755 ;
    END
  END rd_out[158]
  PIN rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.385 0.070 518.455 ;
    END
  END rd_out[159]
  PIN rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.085 0.070 519.155 ;
    END
  END rd_out[160]
  PIN rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.785 0.070 519.855 ;
    END
  END rd_out[161]
  PIN rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.485 0.070 520.555 ;
    END
  END rd_out[162]
  PIN rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.185 0.070 521.255 ;
    END
  END rd_out[163]
  PIN rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.885 0.070 521.955 ;
    END
  END rd_out[164]
  PIN rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.585 0.070 522.655 ;
    END
  END rd_out[165]
  PIN rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.285 0.070 523.355 ;
    END
  END rd_out[166]
  PIN rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.985 0.070 524.055 ;
    END
  END rd_out[167]
  PIN rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.685 0.070 524.755 ;
    END
  END rd_out[168]
  PIN rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.385 0.070 525.455 ;
    END
  END rd_out[169]
  PIN rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.085 0.070 526.155 ;
    END
  END rd_out[170]
  PIN rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.785 0.070 526.855 ;
    END
  END rd_out[171]
  PIN rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.485 0.070 527.555 ;
    END
  END rd_out[172]
  PIN rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.185 0.070 528.255 ;
    END
  END rd_out[173]
  PIN rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.885 0.070 528.955 ;
    END
  END rd_out[174]
  PIN rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.585 0.070 529.655 ;
    END
  END rd_out[175]
  PIN rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.285 0.070 530.355 ;
    END
  END rd_out[176]
  PIN rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.985 0.070 531.055 ;
    END
  END rd_out[177]
  PIN rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.685 0.070 531.755 ;
    END
  END rd_out[178]
  PIN rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.385 0.070 532.455 ;
    END
  END rd_out[179]
  PIN rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.085 0.070 533.155 ;
    END
  END rd_out[180]
  PIN rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.785 0.070 533.855 ;
    END
  END rd_out[181]
  PIN rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.485 0.070 534.555 ;
    END
  END rd_out[182]
  PIN rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.185 0.070 535.255 ;
    END
  END rd_out[183]
  PIN rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.885 0.070 535.955 ;
    END
  END rd_out[184]
  PIN rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.585 0.070 536.655 ;
    END
  END rd_out[185]
  PIN rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.285 0.070 537.355 ;
    END
  END rd_out[186]
  PIN rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.985 0.070 538.055 ;
    END
  END rd_out[187]
  PIN rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.685 0.070 538.755 ;
    END
  END rd_out[188]
  PIN rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.385 0.070 539.455 ;
    END
  END rd_out[189]
  PIN rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.085 0.070 540.155 ;
    END
  END rd_out[190]
  PIN rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.785 0.070 540.855 ;
    END
  END rd_out[191]
  PIN rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.485 0.070 541.555 ;
    END
  END rd_out[192]
  PIN rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.185 0.070 542.255 ;
    END
  END rd_out[193]
  PIN rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.885 0.070 542.955 ;
    END
  END rd_out[194]
  PIN rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.585 0.070 543.655 ;
    END
  END rd_out[195]
  PIN rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.285 0.070 544.355 ;
    END
  END rd_out[196]
  PIN rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.985 0.070 545.055 ;
    END
  END rd_out[197]
  PIN rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.685 0.070 545.755 ;
    END
  END rd_out[198]
  PIN rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.385 0.070 546.455 ;
    END
  END rd_out[199]
  PIN rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.085 0.070 547.155 ;
    END
  END rd_out[200]
  PIN rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.785 0.070 547.855 ;
    END
  END rd_out[201]
  PIN rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.485 0.070 548.555 ;
    END
  END rd_out[202]
  PIN rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.185 0.070 549.255 ;
    END
  END rd_out[203]
  PIN rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.885 0.070 549.955 ;
    END
  END rd_out[204]
  PIN rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.585 0.070 550.655 ;
    END
  END rd_out[205]
  PIN rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.285 0.070 551.355 ;
    END
  END rd_out[206]
  PIN rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.985 0.070 552.055 ;
    END
  END rd_out[207]
  PIN rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.685 0.070 552.755 ;
    END
  END rd_out[208]
  PIN rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.385 0.070 553.455 ;
    END
  END rd_out[209]
  PIN rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.085 0.070 554.155 ;
    END
  END rd_out[210]
  PIN rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.785 0.070 554.855 ;
    END
  END rd_out[211]
  PIN rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.485 0.070 555.555 ;
    END
  END rd_out[212]
  PIN rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.185 0.070 556.255 ;
    END
  END rd_out[213]
  PIN rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.885 0.070 556.955 ;
    END
  END rd_out[214]
  PIN rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.585 0.070 557.655 ;
    END
  END rd_out[215]
  PIN rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.285 0.070 558.355 ;
    END
  END rd_out[216]
  PIN rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.985 0.070 559.055 ;
    END
  END rd_out[217]
  PIN rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.685 0.070 559.755 ;
    END
  END rd_out[218]
  PIN rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.385 0.070 560.455 ;
    END
  END rd_out[219]
  PIN rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.085 0.070 561.155 ;
    END
  END rd_out[220]
  PIN rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.785 0.070 561.855 ;
    END
  END rd_out[221]
  PIN rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.485 0.070 562.555 ;
    END
  END rd_out[222]
  PIN rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.185 0.070 563.255 ;
    END
  END rd_out[223]
  PIN rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.885 0.070 563.955 ;
    END
  END rd_out[224]
  PIN rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.585 0.070 564.655 ;
    END
  END rd_out[225]
  PIN rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.285 0.070 565.355 ;
    END
  END rd_out[226]
  PIN rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.985 0.070 566.055 ;
    END
  END rd_out[227]
  PIN rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.685 0.070 566.755 ;
    END
  END rd_out[228]
  PIN rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.385 0.070 567.455 ;
    END
  END rd_out[229]
  PIN rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.085 0.070 568.155 ;
    END
  END rd_out[230]
  PIN rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.785 0.070 568.855 ;
    END
  END rd_out[231]
  PIN rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.485 0.070 569.555 ;
    END
  END rd_out[232]
  PIN rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.185 0.070 570.255 ;
    END
  END rd_out[233]
  PIN rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.885 0.070 570.955 ;
    END
  END rd_out[234]
  PIN rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.585 0.070 571.655 ;
    END
  END rd_out[235]
  PIN rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.285 0.070 572.355 ;
    END
  END rd_out[236]
  PIN rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.985 0.070 573.055 ;
    END
  END rd_out[237]
  PIN rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.685 0.070 573.755 ;
    END
  END rd_out[238]
  PIN rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.385 0.070 574.455 ;
    END
  END rd_out[239]
  PIN rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.085 0.070 575.155 ;
    END
  END rd_out[240]
  PIN rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.785 0.070 575.855 ;
    END
  END rd_out[241]
  PIN rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.485 0.070 576.555 ;
    END
  END rd_out[242]
  PIN rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.185 0.070 577.255 ;
    END
  END rd_out[243]
  PIN rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.885 0.070 577.955 ;
    END
  END rd_out[244]
  PIN rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.585 0.070 578.655 ;
    END
  END rd_out[245]
  PIN rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.285 0.070 579.355 ;
    END
  END rd_out[246]
  PIN rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.985 0.070 580.055 ;
    END
  END rd_out[247]
  PIN rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.685 0.070 580.755 ;
    END
  END rd_out[248]
  PIN rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.385 0.070 581.455 ;
    END
  END rd_out[249]
  PIN rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.085 0.070 582.155 ;
    END
  END rd_out[250]
  PIN rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.785 0.070 582.855 ;
    END
  END rd_out[251]
  PIN rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.485 0.070 583.555 ;
    END
  END rd_out[252]
  PIN rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.185 0.070 584.255 ;
    END
  END rd_out[253]
  PIN rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.885 0.070 584.955 ;
    END
  END rd_out[254]
  PIN rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.585 0.070 585.655 ;
    END
  END rd_out[255]
  PIN rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.285 0.070 586.355 ;
    END
  END rd_out[256]
  PIN rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.985 0.070 587.055 ;
    END
  END rd_out[257]
  PIN rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.685 0.070 587.755 ;
    END
  END rd_out[258]
  PIN rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.385 0.070 588.455 ;
    END
  END rd_out[259]
  PIN rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.085 0.070 589.155 ;
    END
  END rd_out[260]
  PIN rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.785 0.070 589.855 ;
    END
  END rd_out[261]
  PIN rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.485 0.070 590.555 ;
    END
  END rd_out[262]
  PIN rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.185 0.070 591.255 ;
    END
  END rd_out[263]
  PIN rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.885 0.070 591.955 ;
    END
  END rd_out[264]
  PIN rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.585 0.070 592.655 ;
    END
  END rd_out[265]
  PIN rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.285 0.070 593.355 ;
    END
  END rd_out[266]
  PIN rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.985 0.070 594.055 ;
    END
  END rd_out[267]
  PIN rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.685 0.070 594.755 ;
    END
  END rd_out[268]
  PIN rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.385 0.070 595.455 ;
    END
  END rd_out[269]
  PIN rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.085 0.070 596.155 ;
    END
  END rd_out[270]
  PIN rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.785 0.070 596.855 ;
    END
  END rd_out[271]
  PIN rd_out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.485 0.070 597.555 ;
    END
  END rd_out[272]
  PIN rd_out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.185 0.070 598.255 ;
    END
  END rd_out[273]
  PIN rd_out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.885 0.070 598.955 ;
    END
  END rd_out[274]
  PIN rd_out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.585 0.070 599.655 ;
    END
  END rd_out[275]
  PIN rd_out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.285 0.070 600.355 ;
    END
  END rd_out[276]
  PIN rd_out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.985 0.070 601.055 ;
    END
  END rd_out[277]
  PIN rd_out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.685 0.070 601.755 ;
    END
  END rd_out[278]
  PIN rd_out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.385 0.070 602.455 ;
    END
  END rd_out[279]
  PIN rd_out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.085 0.070 603.155 ;
    END
  END rd_out[280]
  PIN rd_out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.785 0.070 603.855 ;
    END
  END rd_out[281]
  PIN rd_out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.485 0.070 604.555 ;
    END
  END rd_out[282]
  PIN rd_out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.185 0.070 605.255 ;
    END
  END rd_out[283]
  PIN rd_out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.885 0.070 605.955 ;
    END
  END rd_out[284]
  PIN rd_out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.585 0.070 606.655 ;
    END
  END rd_out[285]
  PIN rd_out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.285 0.070 607.355 ;
    END
  END rd_out[286]
  PIN rd_out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.985 0.070 608.055 ;
    END
  END rd_out[287]
  PIN rd_out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.685 0.070 608.755 ;
    END
  END rd_out[288]
  PIN rd_out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.385 0.070 609.455 ;
    END
  END rd_out[289]
  PIN rd_out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.085 0.070 610.155 ;
    END
  END rd_out[290]
  PIN rd_out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.785 0.070 610.855 ;
    END
  END rd_out[291]
  PIN rd_out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.485 0.070 611.555 ;
    END
  END rd_out[292]
  PIN rd_out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.185 0.070 612.255 ;
    END
  END rd_out[293]
  PIN rd_out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.885 0.070 612.955 ;
    END
  END rd_out[294]
  PIN rd_out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.585 0.070 613.655 ;
    END
  END rd_out[295]
  PIN rd_out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.285 0.070 614.355 ;
    END
  END rd_out[296]
  PIN rd_out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.985 0.070 615.055 ;
    END
  END rd_out[297]
  PIN rd_out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.685 0.070 615.755 ;
    END
  END rd_out[298]
  PIN rd_out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.385 0.070 616.455 ;
    END
  END rd_out[299]
  PIN rd_out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.085 0.070 617.155 ;
    END
  END rd_out[300]
  PIN rd_out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.785 0.070 617.855 ;
    END
  END rd_out[301]
  PIN rd_out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.485 0.070 618.555 ;
    END
  END rd_out[302]
  PIN rd_out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.185 0.070 619.255 ;
    END
  END rd_out[303]
  PIN rd_out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.885 0.070 619.955 ;
    END
  END rd_out[304]
  PIN rd_out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.585 0.070 620.655 ;
    END
  END rd_out[305]
  PIN rd_out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.285 0.070 621.355 ;
    END
  END rd_out[306]
  PIN rd_out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.985 0.070 622.055 ;
    END
  END rd_out[307]
  PIN rd_out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.685 0.070 622.755 ;
    END
  END rd_out[308]
  PIN rd_out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.385 0.070 623.455 ;
    END
  END rd_out[309]
  PIN rd_out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.085 0.070 624.155 ;
    END
  END rd_out[310]
  PIN rd_out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.785 0.070 624.855 ;
    END
  END rd_out[311]
  PIN rd_out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.485 0.070 625.555 ;
    END
  END rd_out[312]
  PIN rd_out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.185 0.070 626.255 ;
    END
  END rd_out[313]
  PIN rd_out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.885 0.070 626.955 ;
    END
  END rd_out[314]
  PIN rd_out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.585 0.070 627.655 ;
    END
  END rd_out[315]
  PIN rd_out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.285 0.070 628.355 ;
    END
  END rd_out[316]
  PIN rd_out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.985 0.070 629.055 ;
    END
  END rd_out[317]
  PIN rd_out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.685 0.070 629.755 ;
    END
  END rd_out[318]
  PIN rd_out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.385 0.070 630.455 ;
    END
  END rd_out[319]
  PIN rd_out[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.085 0.070 631.155 ;
    END
  END rd_out[320]
  PIN rd_out[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.785 0.070 631.855 ;
    END
  END rd_out[321]
  PIN rd_out[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.485 0.070 632.555 ;
    END
  END rd_out[322]
  PIN rd_out[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.185 0.070 633.255 ;
    END
  END rd_out[323]
  PIN rd_out[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.885 0.070 633.955 ;
    END
  END rd_out[324]
  PIN rd_out[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.585 0.070 634.655 ;
    END
  END rd_out[325]
  PIN rd_out[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.285 0.070 635.355 ;
    END
  END rd_out[326]
  PIN rd_out[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.985 0.070 636.055 ;
    END
  END rd_out[327]
  PIN rd_out[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.685 0.070 636.755 ;
    END
  END rd_out[328]
  PIN rd_out[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.385 0.070 637.455 ;
    END
  END rd_out[329]
  PIN rd_out[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.085 0.070 638.155 ;
    END
  END rd_out[330]
  PIN rd_out[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.785 0.070 638.855 ;
    END
  END rd_out[331]
  PIN rd_out[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.485 0.070 639.555 ;
    END
  END rd_out[332]
  PIN rd_out[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.185 0.070 640.255 ;
    END
  END rd_out[333]
  PIN rd_out[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.885 0.070 640.955 ;
    END
  END rd_out[334]
  PIN rd_out[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.585 0.070 641.655 ;
    END
  END rd_out[335]
  PIN rd_out[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.285 0.070 642.355 ;
    END
  END rd_out[336]
  PIN rd_out[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.985 0.070 643.055 ;
    END
  END rd_out[337]
  PIN rd_out[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.685 0.070 643.755 ;
    END
  END rd_out[338]
  PIN rd_out[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.385 0.070 644.455 ;
    END
  END rd_out[339]
  PIN rd_out[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.085 0.070 645.155 ;
    END
  END rd_out[340]
  PIN rd_out[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.785 0.070 645.855 ;
    END
  END rd_out[341]
  PIN rd_out[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.485 0.070 646.555 ;
    END
  END rd_out[342]
  PIN rd_out[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.185 0.070 647.255 ;
    END
  END rd_out[343]
  PIN rd_out[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.885 0.070 647.955 ;
    END
  END rd_out[344]
  PIN rd_out[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.585 0.070 648.655 ;
    END
  END rd_out[345]
  PIN rd_out[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.285 0.070 649.355 ;
    END
  END rd_out[346]
  PIN rd_out[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.985 0.070 650.055 ;
    END
  END rd_out[347]
  PIN rd_out[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.685 0.070 650.755 ;
    END
  END rd_out[348]
  PIN rd_out[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.385 0.070 651.455 ;
    END
  END rd_out[349]
  PIN rd_out[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.085 0.070 652.155 ;
    END
  END rd_out[350]
  PIN rd_out[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.785 0.070 652.855 ;
    END
  END rd_out[351]
  PIN rd_out[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.485 0.070 653.555 ;
    END
  END rd_out[352]
  PIN rd_out[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.185 0.070 654.255 ;
    END
  END rd_out[353]
  PIN rd_out[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.885 0.070 654.955 ;
    END
  END rd_out[354]
  PIN rd_out[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.585 0.070 655.655 ;
    END
  END rd_out[355]
  PIN rd_out[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.285 0.070 656.355 ;
    END
  END rd_out[356]
  PIN rd_out[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.985 0.070 657.055 ;
    END
  END rd_out[357]
  PIN rd_out[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.685 0.070 657.755 ;
    END
  END rd_out[358]
  PIN rd_out[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.385 0.070 658.455 ;
    END
  END rd_out[359]
  PIN rd_out[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.085 0.070 659.155 ;
    END
  END rd_out[360]
  PIN rd_out[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.785 0.070 659.855 ;
    END
  END rd_out[361]
  PIN rd_out[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.485 0.070 660.555 ;
    END
  END rd_out[362]
  PIN rd_out[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.185 0.070 661.255 ;
    END
  END rd_out[363]
  PIN rd_out[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.885 0.070 661.955 ;
    END
  END rd_out[364]
  PIN rd_out[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.585 0.070 662.655 ;
    END
  END rd_out[365]
  PIN rd_out[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.285 0.070 663.355 ;
    END
  END rd_out[366]
  PIN rd_out[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.985 0.070 664.055 ;
    END
  END rd_out[367]
  PIN rd_out[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.685 0.070 664.755 ;
    END
  END rd_out[368]
  PIN rd_out[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.385 0.070 665.455 ;
    END
  END rd_out[369]
  PIN rd_out[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.085 0.070 666.155 ;
    END
  END rd_out[370]
  PIN rd_out[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.785 0.070 666.855 ;
    END
  END rd_out[371]
  PIN rd_out[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.485 0.070 667.555 ;
    END
  END rd_out[372]
  PIN rd_out[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.185 0.070 668.255 ;
    END
  END rd_out[373]
  PIN rd_out[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.885 0.070 668.955 ;
    END
  END rd_out[374]
  PIN rd_out[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.585 0.070 669.655 ;
    END
  END rd_out[375]
  PIN rd_out[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.285 0.070 670.355 ;
    END
  END rd_out[376]
  PIN rd_out[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.985 0.070 671.055 ;
    END
  END rd_out[377]
  PIN rd_out[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.685 0.070 671.755 ;
    END
  END rd_out[378]
  PIN rd_out[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.385 0.070 672.455 ;
    END
  END rd_out[379]
  PIN rd_out[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.085 0.070 673.155 ;
    END
  END rd_out[380]
  PIN rd_out[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.785 0.070 673.855 ;
    END
  END rd_out[381]
  PIN rd_out[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.485 0.070 674.555 ;
    END
  END rd_out[382]
  PIN rd_out[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.185 0.070 675.255 ;
    END
  END rd_out[383]
  PIN rd_out[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.885 0.070 675.955 ;
    END
  END rd_out[384]
  PIN rd_out[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.585 0.070 676.655 ;
    END
  END rd_out[385]
  PIN rd_out[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.285 0.070 677.355 ;
    END
  END rd_out[386]
  PIN rd_out[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.985 0.070 678.055 ;
    END
  END rd_out[387]
  PIN rd_out[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.685 0.070 678.755 ;
    END
  END rd_out[388]
  PIN rd_out[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.385 0.070 679.455 ;
    END
  END rd_out[389]
  PIN rd_out[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.085 0.070 680.155 ;
    END
  END rd_out[390]
  PIN rd_out[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.785 0.070 680.855 ;
    END
  END rd_out[391]
  PIN rd_out[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.485 0.070 681.555 ;
    END
  END rd_out[392]
  PIN rd_out[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.185 0.070 682.255 ;
    END
  END rd_out[393]
  PIN rd_out[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.885 0.070 682.955 ;
    END
  END rd_out[394]
  PIN rd_out[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.585 0.070 683.655 ;
    END
  END rd_out[395]
  PIN rd_out[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.285 0.070 684.355 ;
    END
  END rd_out[396]
  PIN rd_out[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.985 0.070 685.055 ;
    END
  END rd_out[397]
  PIN rd_out[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.685 0.070 685.755 ;
    END
  END rd_out[398]
  PIN rd_out[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.385 0.070 686.455 ;
    END
  END rd_out[399]
  PIN rd_out[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.085 0.070 687.155 ;
    END
  END rd_out[400]
  PIN rd_out[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.785 0.070 687.855 ;
    END
  END rd_out[401]
  PIN rd_out[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.485 0.070 688.555 ;
    END
  END rd_out[402]
  PIN rd_out[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.185 0.070 689.255 ;
    END
  END rd_out[403]
  PIN rd_out[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.885 0.070 689.955 ;
    END
  END rd_out[404]
  PIN rd_out[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.585 0.070 690.655 ;
    END
  END rd_out[405]
  PIN rd_out[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.285 0.070 691.355 ;
    END
  END rd_out[406]
  PIN rd_out[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.985 0.070 692.055 ;
    END
  END rd_out[407]
  PIN rd_out[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.685 0.070 692.755 ;
    END
  END rd_out[408]
  PIN rd_out[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.385 0.070 693.455 ;
    END
  END rd_out[409]
  PIN rd_out[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.085 0.070 694.155 ;
    END
  END rd_out[410]
  PIN rd_out[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.785 0.070 694.855 ;
    END
  END rd_out[411]
  PIN rd_out[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.485 0.070 695.555 ;
    END
  END rd_out[412]
  PIN rd_out[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.185 0.070 696.255 ;
    END
  END rd_out[413]
  PIN rd_out[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.885 0.070 696.955 ;
    END
  END rd_out[414]
  PIN rd_out[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.585 0.070 697.655 ;
    END
  END rd_out[415]
  PIN rd_out[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.285 0.070 698.355 ;
    END
  END rd_out[416]
  PIN rd_out[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.985 0.070 699.055 ;
    END
  END rd_out[417]
  PIN rd_out[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.685 0.070 699.755 ;
    END
  END rd_out[418]
  PIN rd_out[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.385 0.070 700.455 ;
    END
  END rd_out[419]
  PIN rd_out[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.085 0.070 701.155 ;
    END
  END rd_out[420]
  PIN rd_out[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.785 0.070 701.855 ;
    END
  END rd_out[421]
  PIN rd_out[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.485 0.070 702.555 ;
    END
  END rd_out[422]
  PIN rd_out[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.185 0.070 703.255 ;
    END
  END rd_out[423]
  PIN rd_out[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.885 0.070 703.955 ;
    END
  END rd_out[424]
  PIN rd_out[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.585 0.070 704.655 ;
    END
  END rd_out[425]
  PIN rd_out[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.285 0.070 705.355 ;
    END
  END rd_out[426]
  PIN rd_out[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.985 0.070 706.055 ;
    END
  END rd_out[427]
  PIN rd_out[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.685 0.070 706.755 ;
    END
  END rd_out[428]
  PIN rd_out[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.385 0.070 707.455 ;
    END
  END rd_out[429]
  PIN rd_out[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.085 0.070 708.155 ;
    END
  END rd_out[430]
  PIN rd_out[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.785 0.070 708.855 ;
    END
  END rd_out[431]
  PIN rd_out[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.485 0.070 709.555 ;
    END
  END rd_out[432]
  PIN rd_out[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.185 0.070 710.255 ;
    END
  END rd_out[433]
  PIN rd_out[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.885 0.070 710.955 ;
    END
  END rd_out[434]
  PIN rd_out[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.585 0.070 711.655 ;
    END
  END rd_out[435]
  PIN rd_out[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.285 0.070 712.355 ;
    END
  END rd_out[436]
  PIN rd_out[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.985 0.070 713.055 ;
    END
  END rd_out[437]
  PIN rd_out[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.685 0.070 713.755 ;
    END
  END rd_out[438]
  PIN rd_out[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.385 0.070 714.455 ;
    END
  END rd_out[439]
  PIN rd_out[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.085 0.070 715.155 ;
    END
  END rd_out[440]
  PIN rd_out[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.785 0.070 715.855 ;
    END
  END rd_out[441]
  PIN rd_out[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.485 0.070 716.555 ;
    END
  END rd_out[442]
  PIN rd_out[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.185 0.070 717.255 ;
    END
  END rd_out[443]
  PIN rd_out[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.885 0.070 717.955 ;
    END
  END rd_out[444]
  PIN rd_out[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.585 0.070 718.655 ;
    END
  END rd_out[445]
  PIN rd_out[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.285 0.070 719.355 ;
    END
  END rd_out[446]
  PIN rd_out[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.985 0.070 720.055 ;
    END
  END rd_out[447]
  PIN rd_out[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.685 0.070 720.755 ;
    END
  END rd_out[448]
  PIN rd_out[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.385 0.070 721.455 ;
    END
  END rd_out[449]
  PIN rd_out[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.085 0.070 722.155 ;
    END
  END rd_out[450]
  PIN rd_out[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.785 0.070 722.855 ;
    END
  END rd_out[451]
  PIN rd_out[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.485 0.070 723.555 ;
    END
  END rd_out[452]
  PIN rd_out[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.185 0.070 724.255 ;
    END
  END rd_out[453]
  PIN rd_out[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.885 0.070 724.955 ;
    END
  END rd_out[454]
  PIN rd_out[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.585 0.070 725.655 ;
    END
  END rd_out[455]
  PIN rd_out[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.285 0.070 726.355 ;
    END
  END rd_out[456]
  PIN rd_out[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.985 0.070 727.055 ;
    END
  END rd_out[457]
  PIN rd_out[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.685 0.070 727.755 ;
    END
  END rd_out[458]
  PIN rd_out[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.385 0.070 728.455 ;
    END
  END rd_out[459]
  PIN rd_out[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.085 0.070 729.155 ;
    END
  END rd_out[460]
  PIN rd_out[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.785 0.070 729.855 ;
    END
  END rd_out[461]
  PIN rd_out[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.485 0.070 730.555 ;
    END
  END rd_out[462]
  PIN rd_out[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.185 0.070 731.255 ;
    END
  END rd_out[463]
  PIN rd_out[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.885 0.070 731.955 ;
    END
  END rd_out[464]
  PIN rd_out[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.585 0.070 732.655 ;
    END
  END rd_out[465]
  PIN rd_out[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.285 0.070 733.355 ;
    END
  END rd_out[466]
  PIN rd_out[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.985 0.070 734.055 ;
    END
  END rd_out[467]
  PIN rd_out[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.685 0.070 734.755 ;
    END
  END rd_out[468]
  PIN rd_out[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.385 0.070 735.455 ;
    END
  END rd_out[469]
  PIN rd_out[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.085 0.070 736.155 ;
    END
  END rd_out[470]
  PIN rd_out[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.785 0.070 736.855 ;
    END
  END rd_out[471]
  PIN rd_out[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.485 0.070 737.555 ;
    END
  END rd_out[472]
  PIN rd_out[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.185 0.070 738.255 ;
    END
  END rd_out[473]
  PIN rd_out[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.885 0.070 738.955 ;
    END
  END rd_out[474]
  PIN rd_out[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.585 0.070 739.655 ;
    END
  END rd_out[475]
  PIN rd_out[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.285 0.070 740.355 ;
    END
  END rd_out[476]
  PIN rd_out[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.985 0.070 741.055 ;
    END
  END rd_out[477]
  PIN rd_out[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.685 0.070 741.755 ;
    END
  END rd_out[478]
  PIN rd_out[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.385 0.070 742.455 ;
    END
  END rd_out[479]
  PIN rd_out[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.085 0.070 743.155 ;
    END
  END rd_out[480]
  PIN rd_out[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.785 0.070 743.855 ;
    END
  END rd_out[481]
  PIN rd_out[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.485 0.070 744.555 ;
    END
  END rd_out[482]
  PIN rd_out[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.185 0.070 745.255 ;
    END
  END rd_out[483]
  PIN rd_out[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.885 0.070 745.955 ;
    END
  END rd_out[484]
  PIN rd_out[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.585 0.070 746.655 ;
    END
  END rd_out[485]
  PIN rd_out[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.285 0.070 747.355 ;
    END
  END rd_out[486]
  PIN rd_out[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.985 0.070 748.055 ;
    END
  END rd_out[487]
  PIN rd_out[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.685 0.070 748.755 ;
    END
  END rd_out[488]
  PIN rd_out[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.385 0.070 749.455 ;
    END
  END rd_out[489]
  PIN rd_out[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.085 0.070 750.155 ;
    END
  END rd_out[490]
  PIN rd_out[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.785 0.070 750.855 ;
    END
  END rd_out[491]
  PIN rd_out[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.485 0.070 751.555 ;
    END
  END rd_out[492]
  PIN rd_out[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.185 0.070 752.255 ;
    END
  END rd_out[493]
  PIN rd_out[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.885 0.070 752.955 ;
    END
  END rd_out[494]
  PIN rd_out[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.585 0.070 753.655 ;
    END
  END rd_out[495]
  PIN rd_out[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.285 0.070 754.355 ;
    END
  END rd_out[496]
  PIN rd_out[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.985 0.070 755.055 ;
    END
  END rd_out[497]
  PIN rd_out[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.685 0.070 755.755 ;
    END
  END rd_out[498]
  PIN rd_out[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.385 0.070 756.455 ;
    END
  END rd_out[499]
  PIN rd_out[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.085 0.070 757.155 ;
    END
  END rd_out[500]
  PIN rd_out[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.785 0.070 757.855 ;
    END
  END rd_out[501]
  PIN rd_out[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.485 0.070 758.555 ;
    END
  END rd_out[502]
  PIN rd_out[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.185 0.070 759.255 ;
    END
  END rd_out[503]
  PIN rd_out[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.885 0.070 759.955 ;
    END
  END rd_out[504]
  PIN rd_out[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.585 0.070 760.655 ;
    END
  END rd_out[505]
  PIN rd_out[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.285 0.070 761.355 ;
    END
  END rd_out[506]
  PIN rd_out[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.985 0.070 762.055 ;
    END
  END rd_out[507]
  PIN rd_out[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.685 0.070 762.755 ;
    END
  END rd_out[508]
  PIN rd_out[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.385 0.070 763.455 ;
    END
  END rd_out[509]
  PIN rd_out[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.085 0.070 764.155 ;
    END
  END rd_out[510]
  PIN rd_out[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.785 0.070 764.855 ;
    END
  END rd_out[511]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.805 0.070 812.875 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.505 0.070 813.575 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.205 0.070 814.275 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.905 0.070 814.975 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.605 0.070 815.675 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.305 0.070 816.375 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.005 0.070 817.075 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.705 0.070 817.775 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.405 0.070 818.475 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.105 0.070 819.175 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.805 0.070 819.875 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.505 0.070 820.575 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.205 0.070 821.275 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.905 0.070 821.975 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.605 0.070 822.675 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.305 0.070 823.375 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.005 0.070 824.075 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.705 0.070 824.775 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.405 0.070 825.475 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.105 0.070 826.175 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.805 0.070 826.875 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.505 0.070 827.575 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.205 0.070 828.275 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.905 0.070 828.975 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.605 0.070 829.675 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.305 0.070 830.375 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.005 0.070 831.075 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.705 0.070 831.775 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.405 0.070 832.475 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.105 0.070 833.175 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.805 0.070 833.875 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.505 0.070 834.575 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.205 0.070 835.275 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.905 0.070 835.975 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.605 0.070 836.675 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.305 0.070 837.375 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.005 0.070 838.075 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.705 0.070 838.775 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.405 0.070 839.475 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.105 0.070 840.175 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.805 0.070 840.875 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.505 0.070 841.575 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.205 0.070 842.275 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.905 0.070 842.975 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.605 0.070 843.675 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.305 0.070 844.375 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.005 0.070 845.075 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.705 0.070 845.775 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.405 0.070 846.475 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.105 0.070 847.175 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.805 0.070 847.875 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.505 0.070 848.575 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.205 0.070 849.275 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.905 0.070 849.975 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.605 0.070 850.675 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.305 0.070 851.375 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.005 0.070 852.075 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.705 0.070 852.775 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.405 0.070 853.475 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.105 0.070 854.175 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.805 0.070 854.875 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.505 0.070 855.575 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.205 0.070 856.275 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.905 0.070 856.975 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.605 0.070 857.675 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.305 0.070 858.375 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.005 0.070 859.075 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.705 0.070 859.775 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.405 0.070 860.475 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.105 0.070 861.175 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.805 0.070 861.875 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.505 0.070 862.575 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.205 0.070 863.275 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.905 0.070 863.975 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.605 0.070 864.675 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.305 0.070 865.375 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.005 0.070 866.075 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.705 0.070 866.775 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.405 0.070 867.475 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.105 0.070 868.175 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.805 0.070 868.875 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.505 0.070 869.575 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.205 0.070 870.275 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.905 0.070 870.975 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.605 0.070 871.675 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.305 0.070 872.375 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.005 0.070 873.075 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.705 0.070 873.775 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.405 0.070 874.475 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.105 0.070 875.175 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.805 0.070 875.875 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.505 0.070 876.575 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.205 0.070 877.275 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.905 0.070 877.975 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.605 0.070 878.675 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.305 0.070 879.375 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.005 0.070 880.075 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.705 0.070 880.775 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.405 0.070 881.475 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.105 0.070 882.175 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.805 0.070 882.875 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.505 0.070 883.575 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.205 0.070 884.275 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.905 0.070 884.975 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.605 0.070 885.675 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.305 0.070 886.375 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.005 0.070 887.075 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.705 0.070 887.775 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.405 0.070 888.475 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.105 0.070 889.175 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.805 0.070 889.875 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.505 0.070 890.575 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.205 0.070 891.275 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.905 0.070 891.975 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.605 0.070 892.675 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.305 0.070 893.375 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.005 0.070 894.075 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.705 0.070 894.775 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.405 0.070 895.475 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.105 0.070 896.175 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.805 0.070 896.875 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.505 0.070 897.575 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.205 0.070 898.275 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.905 0.070 898.975 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.605 0.070 899.675 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.305 0.070 900.375 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.005 0.070 901.075 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.705 0.070 901.775 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.405 0.070 902.475 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 903.105 0.070 903.175 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 903.805 0.070 903.875 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 904.505 0.070 904.575 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 905.205 0.070 905.275 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 905.905 0.070 905.975 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 906.605 0.070 906.675 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 907.305 0.070 907.375 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 908.005 0.070 908.075 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 908.705 0.070 908.775 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 909.405 0.070 909.475 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 910.105 0.070 910.175 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 910.805 0.070 910.875 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 911.505 0.070 911.575 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 912.205 0.070 912.275 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 912.905 0.070 912.975 ;
    END
  END wd_in[143]
  PIN wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 913.605 0.070 913.675 ;
    END
  END wd_in[144]
  PIN wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 914.305 0.070 914.375 ;
    END
  END wd_in[145]
  PIN wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 915.005 0.070 915.075 ;
    END
  END wd_in[146]
  PIN wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 915.705 0.070 915.775 ;
    END
  END wd_in[147]
  PIN wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 916.405 0.070 916.475 ;
    END
  END wd_in[148]
  PIN wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 917.105 0.070 917.175 ;
    END
  END wd_in[149]
  PIN wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 917.805 0.070 917.875 ;
    END
  END wd_in[150]
  PIN wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 918.505 0.070 918.575 ;
    END
  END wd_in[151]
  PIN wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 919.205 0.070 919.275 ;
    END
  END wd_in[152]
  PIN wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 919.905 0.070 919.975 ;
    END
  END wd_in[153]
  PIN wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 920.605 0.070 920.675 ;
    END
  END wd_in[154]
  PIN wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 921.305 0.070 921.375 ;
    END
  END wd_in[155]
  PIN wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 922.005 0.070 922.075 ;
    END
  END wd_in[156]
  PIN wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 922.705 0.070 922.775 ;
    END
  END wd_in[157]
  PIN wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 923.405 0.070 923.475 ;
    END
  END wd_in[158]
  PIN wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 924.105 0.070 924.175 ;
    END
  END wd_in[159]
  PIN wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 924.805 0.070 924.875 ;
    END
  END wd_in[160]
  PIN wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 925.505 0.070 925.575 ;
    END
  END wd_in[161]
  PIN wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 926.205 0.070 926.275 ;
    END
  END wd_in[162]
  PIN wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 926.905 0.070 926.975 ;
    END
  END wd_in[163]
  PIN wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 927.605 0.070 927.675 ;
    END
  END wd_in[164]
  PIN wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 928.305 0.070 928.375 ;
    END
  END wd_in[165]
  PIN wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 929.005 0.070 929.075 ;
    END
  END wd_in[166]
  PIN wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 929.705 0.070 929.775 ;
    END
  END wd_in[167]
  PIN wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 930.405 0.070 930.475 ;
    END
  END wd_in[168]
  PIN wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 931.105 0.070 931.175 ;
    END
  END wd_in[169]
  PIN wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 931.805 0.070 931.875 ;
    END
  END wd_in[170]
  PIN wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 932.505 0.070 932.575 ;
    END
  END wd_in[171]
  PIN wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 933.205 0.070 933.275 ;
    END
  END wd_in[172]
  PIN wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 933.905 0.070 933.975 ;
    END
  END wd_in[173]
  PIN wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 934.605 0.070 934.675 ;
    END
  END wd_in[174]
  PIN wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 935.305 0.070 935.375 ;
    END
  END wd_in[175]
  PIN wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 936.005 0.070 936.075 ;
    END
  END wd_in[176]
  PIN wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 936.705 0.070 936.775 ;
    END
  END wd_in[177]
  PIN wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 937.405 0.070 937.475 ;
    END
  END wd_in[178]
  PIN wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 938.105 0.070 938.175 ;
    END
  END wd_in[179]
  PIN wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 938.805 0.070 938.875 ;
    END
  END wd_in[180]
  PIN wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 939.505 0.070 939.575 ;
    END
  END wd_in[181]
  PIN wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 940.205 0.070 940.275 ;
    END
  END wd_in[182]
  PIN wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 940.905 0.070 940.975 ;
    END
  END wd_in[183]
  PIN wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 941.605 0.070 941.675 ;
    END
  END wd_in[184]
  PIN wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 942.305 0.070 942.375 ;
    END
  END wd_in[185]
  PIN wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 943.005 0.070 943.075 ;
    END
  END wd_in[186]
  PIN wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 943.705 0.070 943.775 ;
    END
  END wd_in[187]
  PIN wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 944.405 0.070 944.475 ;
    END
  END wd_in[188]
  PIN wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 945.105 0.070 945.175 ;
    END
  END wd_in[189]
  PIN wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 945.805 0.070 945.875 ;
    END
  END wd_in[190]
  PIN wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 946.505 0.070 946.575 ;
    END
  END wd_in[191]
  PIN wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 947.205 0.070 947.275 ;
    END
  END wd_in[192]
  PIN wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 947.905 0.070 947.975 ;
    END
  END wd_in[193]
  PIN wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 948.605 0.070 948.675 ;
    END
  END wd_in[194]
  PIN wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 949.305 0.070 949.375 ;
    END
  END wd_in[195]
  PIN wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 950.005 0.070 950.075 ;
    END
  END wd_in[196]
  PIN wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 950.705 0.070 950.775 ;
    END
  END wd_in[197]
  PIN wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 951.405 0.070 951.475 ;
    END
  END wd_in[198]
  PIN wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 952.105 0.070 952.175 ;
    END
  END wd_in[199]
  PIN wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 952.805 0.070 952.875 ;
    END
  END wd_in[200]
  PIN wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 953.505 0.070 953.575 ;
    END
  END wd_in[201]
  PIN wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 954.205 0.070 954.275 ;
    END
  END wd_in[202]
  PIN wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 954.905 0.070 954.975 ;
    END
  END wd_in[203]
  PIN wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 955.605 0.070 955.675 ;
    END
  END wd_in[204]
  PIN wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 956.305 0.070 956.375 ;
    END
  END wd_in[205]
  PIN wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 957.005 0.070 957.075 ;
    END
  END wd_in[206]
  PIN wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 957.705 0.070 957.775 ;
    END
  END wd_in[207]
  PIN wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 958.405 0.070 958.475 ;
    END
  END wd_in[208]
  PIN wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 959.105 0.070 959.175 ;
    END
  END wd_in[209]
  PIN wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 959.805 0.070 959.875 ;
    END
  END wd_in[210]
  PIN wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 960.505 0.070 960.575 ;
    END
  END wd_in[211]
  PIN wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 961.205 0.070 961.275 ;
    END
  END wd_in[212]
  PIN wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 961.905 0.070 961.975 ;
    END
  END wd_in[213]
  PIN wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 962.605 0.070 962.675 ;
    END
  END wd_in[214]
  PIN wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 963.305 0.070 963.375 ;
    END
  END wd_in[215]
  PIN wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 964.005 0.070 964.075 ;
    END
  END wd_in[216]
  PIN wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 964.705 0.070 964.775 ;
    END
  END wd_in[217]
  PIN wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 965.405 0.070 965.475 ;
    END
  END wd_in[218]
  PIN wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 966.105 0.070 966.175 ;
    END
  END wd_in[219]
  PIN wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 966.805 0.070 966.875 ;
    END
  END wd_in[220]
  PIN wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 967.505 0.070 967.575 ;
    END
  END wd_in[221]
  PIN wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 968.205 0.070 968.275 ;
    END
  END wd_in[222]
  PIN wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 968.905 0.070 968.975 ;
    END
  END wd_in[223]
  PIN wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 969.605 0.070 969.675 ;
    END
  END wd_in[224]
  PIN wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 970.305 0.070 970.375 ;
    END
  END wd_in[225]
  PIN wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 971.005 0.070 971.075 ;
    END
  END wd_in[226]
  PIN wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 971.705 0.070 971.775 ;
    END
  END wd_in[227]
  PIN wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 972.405 0.070 972.475 ;
    END
  END wd_in[228]
  PIN wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 973.105 0.070 973.175 ;
    END
  END wd_in[229]
  PIN wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 973.805 0.070 973.875 ;
    END
  END wd_in[230]
  PIN wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 974.505 0.070 974.575 ;
    END
  END wd_in[231]
  PIN wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 975.205 0.070 975.275 ;
    END
  END wd_in[232]
  PIN wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 975.905 0.070 975.975 ;
    END
  END wd_in[233]
  PIN wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 976.605 0.070 976.675 ;
    END
  END wd_in[234]
  PIN wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 977.305 0.070 977.375 ;
    END
  END wd_in[235]
  PIN wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 978.005 0.070 978.075 ;
    END
  END wd_in[236]
  PIN wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 978.705 0.070 978.775 ;
    END
  END wd_in[237]
  PIN wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 979.405 0.070 979.475 ;
    END
  END wd_in[238]
  PIN wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 980.105 0.070 980.175 ;
    END
  END wd_in[239]
  PIN wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 980.805 0.070 980.875 ;
    END
  END wd_in[240]
  PIN wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 981.505 0.070 981.575 ;
    END
  END wd_in[241]
  PIN wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 982.205 0.070 982.275 ;
    END
  END wd_in[242]
  PIN wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 982.905 0.070 982.975 ;
    END
  END wd_in[243]
  PIN wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 983.605 0.070 983.675 ;
    END
  END wd_in[244]
  PIN wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 984.305 0.070 984.375 ;
    END
  END wd_in[245]
  PIN wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 985.005 0.070 985.075 ;
    END
  END wd_in[246]
  PIN wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 985.705 0.070 985.775 ;
    END
  END wd_in[247]
  PIN wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 986.405 0.070 986.475 ;
    END
  END wd_in[248]
  PIN wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 987.105 0.070 987.175 ;
    END
  END wd_in[249]
  PIN wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 987.805 0.070 987.875 ;
    END
  END wd_in[250]
  PIN wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 988.505 0.070 988.575 ;
    END
  END wd_in[251]
  PIN wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 989.205 0.070 989.275 ;
    END
  END wd_in[252]
  PIN wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 989.905 0.070 989.975 ;
    END
  END wd_in[253]
  PIN wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 990.605 0.070 990.675 ;
    END
  END wd_in[254]
  PIN wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 991.305 0.070 991.375 ;
    END
  END wd_in[255]
  PIN wd_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 992.005 0.070 992.075 ;
    END
  END wd_in[256]
  PIN wd_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 992.705 0.070 992.775 ;
    END
  END wd_in[257]
  PIN wd_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 993.405 0.070 993.475 ;
    END
  END wd_in[258]
  PIN wd_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 994.105 0.070 994.175 ;
    END
  END wd_in[259]
  PIN wd_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 994.805 0.070 994.875 ;
    END
  END wd_in[260]
  PIN wd_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 995.505 0.070 995.575 ;
    END
  END wd_in[261]
  PIN wd_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 996.205 0.070 996.275 ;
    END
  END wd_in[262]
  PIN wd_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 996.905 0.070 996.975 ;
    END
  END wd_in[263]
  PIN wd_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 997.605 0.070 997.675 ;
    END
  END wd_in[264]
  PIN wd_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 998.305 0.070 998.375 ;
    END
  END wd_in[265]
  PIN wd_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 999.005 0.070 999.075 ;
    END
  END wd_in[266]
  PIN wd_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 999.705 0.070 999.775 ;
    END
  END wd_in[267]
  PIN wd_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1000.405 0.070 1000.475 ;
    END
  END wd_in[268]
  PIN wd_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1001.105 0.070 1001.175 ;
    END
  END wd_in[269]
  PIN wd_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1001.805 0.070 1001.875 ;
    END
  END wd_in[270]
  PIN wd_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1002.505 0.070 1002.575 ;
    END
  END wd_in[271]
  PIN wd_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1003.205 0.070 1003.275 ;
    END
  END wd_in[272]
  PIN wd_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1003.905 0.070 1003.975 ;
    END
  END wd_in[273]
  PIN wd_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1004.605 0.070 1004.675 ;
    END
  END wd_in[274]
  PIN wd_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1005.305 0.070 1005.375 ;
    END
  END wd_in[275]
  PIN wd_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1006.005 0.070 1006.075 ;
    END
  END wd_in[276]
  PIN wd_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1006.705 0.070 1006.775 ;
    END
  END wd_in[277]
  PIN wd_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1007.405 0.070 1007.475 ;
    END
  END wd_in[278]
  PIN wd_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.105 0.070 1008.175 ;
    END
  END wd_in[279]
  PIN wd_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.805 0.070 1008.875 ;
    END
  END wd_in[280]
  PIN wd_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1009.505 0.070 1009.575 ;
    END
  END wd_in[281]
  PIN wd_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.205 0.070 1010.275 ;
    END
  END wd_in[282]
  PIN wd_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.905 0.070 1010.975 ;
    END
  END wd_in[283]
  PIN wd_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1011.605 0.070 1011.675 ;
    END
  END wd_in[284]
  PIN wd_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1012.305 0.070 1012.375 ;
    END
  END wd_in[285]
  PIN wd_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.005 0.070 1013.075 ;
    END
  END wd_in[286]
  PIN wd_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.705 0.070 1013.775 ;
    END
  END wd_in[287]
  PIN wd_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.405 0.070 1014.475 ;
    END
  END wd_in[288]
  PIN wd_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.105 0.070 1015.175 ;
    END
  END wd_in[289]
  PIN wd_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.805 0.070 1015.875 ;
    END
  END wd_in[290]
  PIN wd_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1016.505 0.070 1016.575 ;
    END
  END wd_in[291]
  PIN wd_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.205 0.070 1017.275 ;
    END
  END wd_in[292]
  PIN wd_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.905 0.070 1017.975 ;
    END
  END wd_in[293]
  PIN wd_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1018.605 0.070 1018.675 ;
    END
  END wd_in[294]
  PIN wd_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1019.305 0.070 1019.375 ;
    END
  END wd_in[295]
  PIN wd_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.005 0.070 1020.075 ;
    END
  END wd_in[296]
  PIN wd_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.705 0.070 1020.775 ;
    END
  END wd_in[297]
  PIN wd_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1021.405 0.070 1021.475 ;
    END
  END wd_in[298]
  PIN wd_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.105 0.070 1022.175 ;
    END
  END wd_in[299]
  PIN wd_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.805 0.070 1022.875 ;
    END
  END wd_in[300]
  PIN wd_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1023.505 0.070 1023.575 ;
    END
  END wd_in[301]
  PIN wd_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.205 0.070 1024.275 ;
    END
  END wd_in[302]
  PIN wd_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.905 0.070 1024.975 ;
    END
  END wd_in[303]
  PIN wd_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1025.605 0.070 1025.675 ;
    END
  END wd_in[304]
  PIN wd_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1026.305 0.070 1026.375 ;
    END
  END wd_in[305]
  PIN wd_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.005 0.070 1027.075 ;
    END
  END wd_in[306]
  PIN wd_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.705 0.070 1027.775 ;
    END
  END wd_in[307]
  PIN wd_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1028.405 0.070 1028.475 ;
    END
  END wd_in[308]
  PIN wd_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.105 0.070 1029.175 ;
    END
  END wd_in[309]
  PIN wd_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.805 0.070 1029.875 ;
    END
  END wd_in[310]
  PIN wd_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1030.505 0.070 1030.575 ;
    END
  END wd_in[311]
  PIN wd_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.205 0.070 1031.275 ;
    END
  END wd_in[312]
  PIN wd_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.905 0.070 1031.975 ;
    END
  END wd_in[313]
  PIN wd_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1032.605 0.070 1032.675 ;
    END
  END wd_in[314]
  PIN wd_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1033.305 0.070 1033.375 ;
    END
  END wd_in[315]
  PIN wd_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.005 0.070 1034.075 ;
    END
  END wd_in[316]
  PIN wd_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.705 0.070 1034.775 ;
    END
  END wd_in[317]
  PIN wd_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.405 0.070 1035.475 ;
    END
  END wd_in[318]
  PIN wd_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.105 0.070 1036.175 ;
    END
  END wd_in[319]
  PIN wd_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.805 0.070 1036.875 ;
    END
  END wd_in[320]
  PIN wd_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1037.505 0.070 1037.575 ;
    END
  END wd_in[321]
  PIN wd_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.205 0.070 1038.275 ;
    END
  END wd_in[322]
  PIN wd_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.905 0.070 1038.975 ;
    END
  END wd_in[323]
  PIN wd_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1039.605 0.070 1039.675 ;
    END
  END wd_in[324]
  PIN wd_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1040.305 0.070 1040.375 ;
    END
  END wd_in[325]
  PIN wd_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.005 0.070 1041.075 ;
    END
  END wd_in[326]
  PIN wd_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.705 0.070 1041.775 ;
    END
  END wd_in[327]
  PIN wd_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1042.405 0.070 1042.475 ;
    END
  END wd_in[328]
  PIN wd_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.105 0.070 1043.175 ;
    END
  END wd_in[329]
  PIN wd_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.805 0.070 1043.875 ;
    END
  END wd_in[330]
  PIN wd_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1044.505 0.070 1044.575 ;
    END
  END wd_in[331]
  PIN wd_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.205 0.070 1045.275 ;
    END
  END wd_in[332]
  PIN wd_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.905 0.070 1045.975 ;
    END
  END wd_in[333]
  PIN wd_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.605 0.070 1046.675 ;
    END
  END wd_in[334]
  PIN wd_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1047.305 0.070 1047.375 ;
    END
  END wd_in[335]
  PIN wd_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.005 0.070 1048.075 ;
    END
  END wd_in[336]
  PIN wd_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.705 0.070 1048.775 ;
    END
  END wd_in[337]
  PIN wd_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1049.405 0.070 1049.475 ;
    END
  END wd_in[338]
  PIN wd_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.105 0.070 1050.175 ;
    END
  END wd_in[339]
  PIN wd_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.805 0.070 1050.875 ;
    END
  END wd_in[340]
  PIN wd_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1051.505 0.070 1051.575 ;
    END
  END wd_in[341]
  PIN wd_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.205 0.070 1052.275 ;
    END
  END wd_in[342]
  PIN wd_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.905 0.070 1052.975 ;
    END
  END wd_in[343]
  PIN wd_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1053.605 0.070 1053.675 ;
    END
  END wd_in[344]
  PIN wd_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1054.305 0.070 1054.375 ;
    END
  END wd_in[345]
  PIN wd_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.005 0.070 1055.075 ;
    END
  END wd_in[346]
  PIN wd_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.705 0.070 1055.775 ;
    END
  END wd_in[347]
  PIN wd_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1056.405 0.070 1056.475 ;
    END
  END wd_in[348]
  PIN wd_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.105 0.070 1057.175 ;
    END
  END wd_in[349]
  PIN wd_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.805 0.070 1057.875 ;
    END
  END wd_in[350]
  PIN wd_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1058.505 0.070 1058.575 ;
    END
  END wd_in[351]
  PIN wd_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.205 0.070 1059.275 ;
    END
  END wd_in[352]
  PIN wd_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.905 0.070 1059.975 ;
    END
  END wd_in[353]
  PIN wd_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1060.605 0.070 1060.675 ;
    END
  END wd_in[354]
  PIN wd_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1061.305 0.070 1061.375 ;
    END
  END wd_in[355]
  PIN wd_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.005 0.070 1062.075 ;
    END
  END wd_in[356]
  PIN wd_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.705 0.070 1062.775 ;
    END
  END wd_in[357]
  PIN wd_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1063.405 0.070 1063.475 ;
    END
  END wd_in[358]
  PIN wd_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.105 0.070 1064.175 ;
    END
  END wd_in[359]
  PIN wd_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.805 0.070 1064.875 ;
    END
  END wd_in[360]
  PIN wd_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1065.505 0.070 1065.575 ;
    END
  END wd_in[361]
  PIN wd_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.205 0.070 1066.275 ;
    END
  END wd_in[362]
  PIN wd_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.905 0.070 1066.975 ;
    END
  END wd_in[363]
  PIN wd_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1067.605 0.070 1067.675 ;
    END
  END wd_in[364]
  PIN wd_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.305 0.070 1068.375 ;
    END
  END wd_in[365]
  PIN wd_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.005 0.070 1069.075 ;
    END
  END wd_in[366]
  PIN wd_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.705 0.070 1069.775 ;
    END
  END wd_in[367]
  PIN wd_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1070.405 0.070 1070.475 ;
    END
  END wd_in[368]
  PIN wd_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.105 0.070 1071.175 ;
    END
  END wd_in[369]
  PIN wd_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.805 0.070 1071.875 ;
    END
  END wd_in[370]
  PIN wd_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1072.505 0.070 1072.575 ;
    END
  END wd_in[371]
  PIN wd_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.205 0.070 1073.275 ;
    END
  END wd_in[372]
  PIN wd_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.905 0.070 1073.975 ;
    END
  END wd_in[373]
  PIN wd_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1074.605 0.070 1074.675 ;
    END
  END wd_in[374]
  PIN wd_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1075.305 0.070 1075.375 ;
    END
  END wd_in[375]
  PIN wd_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.005 0.070 1076.075 ;
    END
  END wd_in[376]
  PIN wd_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.705 0.070 1076.775 ;
    END
  END wd_in[377]
  PIN wd_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1077.405 0.070 1077.475 ;
    END
  END wd_in[378]
  PIN wd_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.105 0.070 1078.175 ;
    END
  END wd_in[379]
  PIN wd_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.805 0.070 1078.875 ;
    END
  END wd_in[380]
  PIN wd_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1079.505 0.070 1079.575 ;
    END
  END wd_in[381]
  PIN wd_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.205 0.070 1080.275 ;
    END
  END wd_in[382]
  PIN wd_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.905 0.070 1080.975 ;
    END
  END wd_in[383]
  PIN wd_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1081.605 0.070 1081.675 ;
    END
  END wd_in[384]
  PIN wd_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1082.305 0.070 1082.375 ;
    END
  END wd_in[385]
  PIN wd_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.005 0.070 1083.075 ;
    END
  END wd_in[386]
  PIN wd_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.705 0.070 1083.775 ;
    END
  END wd_in[387]
  PIN wd_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1084.405 0.070 1084.475 ;
    END
  END wd_in[388]
  PIN wd_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.105 0.070 1085.175 ;
    END
  END wd_in[389]
  PIN wd_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.805 0.070 1085.875 ;
    END
  END wd_in[390]
  PIN wd_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1086.505 0.070 1086.575 ;
    END
  END wd_in[391]
  PIN wd_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.205 0.070 1087.275 ;
    END
  END wd_in[392]
  PIN wd_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.905 0.070 1087.975 ;
    END
  END wd_in[393]
  PIN wd_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1088.605 0.070 1088.675 ;
    END
  END wd_in[394]
  PIN wd_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.305 0.070 1089.375 ;
    END
  END wd_in[395]
  PIN wd_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.005 0.070 1090.075 ;
    END
  END wd_in[396]
  PIN wd_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.705 0.070 1090.775 ;
    END
  END wd_in[397]
  PIN wd_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1091.405 0.070 1091.475 ;
    END
  END wd_in[398]
  PIN wd_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.105 0.070 1092.175 ;
    END
  END wd_in[399]
  PIN wd_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.805 0.070 1092.875 ;
    END
  END wd_in[400]
  PIN wd_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1093.505 0.070 1093.575 ;
    END
  END wd_in[401]
  PIN wd_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.205 0.070 1094.275 ;
    END
  END wd_in[402]
  PIN wd_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.905 0.070 1094.975 ;
    END
  END wd_in[403]
  PIN wd_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1095.605 0.070 1095.675 ;
    END
  END wd_in[404]
  PIN wd_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1096.305 0.070 1096.375 ;
    END
  END wd_in[405]
  PIN wd_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.005 0.070 1097.075 ;
    END
  END wd_in[406]
  PIN wd_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.705 0.070 1097.775 ;
    END
  END wd_in[407]
  PIN wd_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1098.405 0.070 1098.475 ;
    END
  END wd_in[408]
  PIN wd_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.105 0.070 1099.175 ;
    END
  END wd_in[409]
  PIN wd_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.805 0.070 1099.875 ;
    END
  END wd_in[410]
  PIN wd_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.505 0.070 1100.575 ;
    END
  END wd_in[411]
  PIN wd_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.205 0.070 1101.275 ;
    END
  END wd_in[412]
  PIN wd_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.905 0.070 1101.975 ;
    END
  END wd_in[413]
  PIN wd_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1102.605 0.070 1102.675 ;
    END
  END wd_in[414]
  PIN wd_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1103.305 0.070 1103.375 ;
    END
  END wd_in[415]
  PIN wd_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.005 0.070 1104.075 ;
    END
  END wd_in[416]
  PIN wd_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.705 0.070 1104.775 ;
    END
  END wd_in[417]
  PIN wd_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1105.405 0.070 1105.475 ;
    END
  END wd_in[418]
  PIN wd_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.105 0.070 1106.175 ;
    END
  END wd_in[419]
  PIN wd_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.805 0.070 1106.875 ;
    END
  END wd_in[420]
  PIN wd_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1107.505 0.070 1107.575 ;
    END
  END wd_in[421]
  PIN wd_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.205 0.070 1108.275 ;
    END
  END wd_in[422]
  PIN wd_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.905 0.070 1108.975 ;
    END
  END wd_in[423]
  PIN wd_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1109.605 0.070 1109.675 ;
    END
  END wd_in[424]
  PIN wd_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1110.305 0.070 1110.375 ;
    END
  END wd_in[425]
  PIN wd_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.005 0.070 1111.075 ;
    END
  END wd_in[426]
  PIN wd_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.705 0.070 1111.775 ;
    END
  END wd_in[427]
  PIN wd_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1112.405 0.070 1112.475 ;
    END
  END wd_in[428]
  PIN wd_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.105 0.070 1113.175 ;
    END
  END wd_in[429]
  PIN wd_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.805 0.070 1113.875 ;
    END
  END wd_in[430]
  PIN wd_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1114.505 0.070 1114.575 ;
    END
  END wd_in[431]
  PIN wd_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.205 0.070 1115.275 ;
    END
  END wd_in[432]
  PIN wd_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.905 0.070 1115.975 ;
    END
  END wd_in[433]
  PIN wd_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1116.605 0.070 1116.675 ;
    END
  END wd_in[434]
  PIN wd_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1117.305 0.070 1117.375 ;
    END
  END wd_in[435]
  PIN wd_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.005 0.070 1118.075 ;
    END
  END wd_in[436]
  PIN wd_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.705 0.070 1118.775 ;
    END
  END wd_in[437]
  PIN wd_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1119.405 0.070 1119.475 ;
    END
  END wd_in[438]
  PIN wd_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.105 0.070 1120.175 ;
    END
  END wd_in[439]
  PIN wd_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.805 0.070 1120.875 ;
    END
  END wd_in[440]
  PIN wd_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.505 0.070 1121.575 ;
    END
  END wd_in[441]
  PIN wd_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.205 0.070 1122.275 ;
    END
  END wd_in[442]
  PIN wd_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.905 0.070 1122.975 ;
    END
  END wd_in[443]
  PIN wd_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1123.605 0.070 1123.675 ;
    END
  END wd_in[444]
  PIN wd_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1124.305 0.070 1124.375 ;
    END
  END wd_in[445]
  PIN wd_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.005 0.070 1125.075 ;
    END
  END wd_in[446]
  PIN wd_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.705 0.070 1125.775 ;
    END
  END wd_in[447]
  PIN wd_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1126.405 0.070 1126.475 ;
    END
  END wd_in[448]
  PIN wd_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.105 0.070 1127.175 ;
    END
  END wd_in[449]
  PIN wd_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.805 0.070 1127.875 ;
    END
  END wd_in[450]
  PIN wd_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1128.505 0.070 1128.575 ;
    END
  END wd_in[451]
  PIN wd_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.205 0.070 1129.275 ;
    END
  END wd_in[452]
  PIN wd_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.905 0.070 1129.975 ;
    END
  END wd_in[453]
  PIN wd_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1130.605 0.070 1130.675 ;
    END
  END wd_in[454]
  PIN wd_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1131.305 0.070 1131.375 ;
    END
  END wd_in[455]
  PIN wd_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.005 0.070 1132.075 ;
    END
  END wd_in[456]
  PIN wd_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.705 0.070 1132.775 ;
    END
  END wd_in[457]
  PIN wd_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1133.405 0.070 1133.475 ;
    END
  END wd_in[458]
  PIN wd_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.105 0.070 1134.175 ;
    END
  END wd_in[459]
  PIN wd_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.805 0.070 1134.875 ;
    END
  END wd_in[460]
  PIN wd_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1135.505 0.070 1135.575 ;
    END
  END wd_in[461]
  PIN wd_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.205 0.070 1136.275 ;
    END
  END wd_in[462]
  PIN wd_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.905 0.070 1136.975 ;
    END
  END wd_in[463]
  PIN wd_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1137.605 0.070 1137.675 ;
    END
  END wd_in[464]
  PIN wd_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1138.305 0.070 1138.375 ;
    END
  END wd_in[465]
  PIN wd_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.005 0.070 1139.075 ;
    END
  END wd_in[466]
  PIN wd_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.705 0.070 1139.775 ;
    END
  END wd_in[467]
  PIN wd_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1140.405 0.070 1140.475 ;
    END
  END wd_in[468]
  PIN wd_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.105 0.070 1141.175 ;
    END
  END wd_in[469]
  PIN wd_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.805 0.070 1141.875 ;
    END
  END wd_in[470]
  PIN wd_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1142.505 0.070 1142.575 ;
    END
  END wd_in[471]
  PIN wd_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.205 0.070 1143.275 ;
    END
  END wd_in[472]
  PIN wd_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.905 0.070 1143.975 ;
    END
  END wd_in[473]
  PIN wd_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1144.605 0.070 1144.675 ;
    END
  END wd_in[474]
  PIN wd_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1145.305 0.070 1145.375 ;
    END
  END wd_in[475]
  PIN wd_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.005 0.070 1146.075 ;
    END
  END wd_in[476]
  PIN wd_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.705 0.070 1146.775 ;
    END
  END wd_in[477]
  PIN wd_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1147.405 0.070 1147.475 ;
    END
  END wd_in[478]
  PIN wd_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.105 0.070 1148.175 ;
    END
  END wd_in[479]
  PIN wd_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.805 0.070 1148.875 ;
    END
  END wd_in[480]
  PIN wd_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1149.505 0.070 1149.575 ;
    END
  END wd_in[481]
  PIN wd_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.205 0.070 1150.275 ;
    END
  END wd_in[482]
  PIN wd_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.905 0.070 1150.975 ;
    END
  END wd_in[483]
  PIN wd_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1151.605 0.070 1151.675 ;
    END
  END wd_in[484]
  PIN wd_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1152.305 0.070 1152.375 ;
    END
  END wd_in[485]
  PIN wd_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.005 0.070 1153.075 ;
    END
  END wd_in[486]
  PIN wd_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.705 0.070 1153.775 ;
    END
  END wd_in[487]
  PIN wd_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.405 0.070 1154.475 ;
    END
  END wd_in[488]
  PIN wd_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.105 0.070 1155.175 ;
    END
  END wd_in[489]
  PIN wd_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.805 0.070 1155.875 ;
    END
  END wd_in[490]
  PIN wd_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1156.505 0.070 1156.575 ;
    END
  END wd_in[491]
  PIN wd_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.205 0.070 1157.275 ;
    END
  END wd_in[492]
  PIN wd_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.905 0.070 1157.975 ;
    END
  END wd_in[493]
  PIN wd_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1158.605 0.070 1158.675 ;
    END
  END wd_in[494]
  PIN wd_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1159.305 0.070 1159.375 ;
    END
  END wd_in[495]
  PIN wd_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.005 0.070 1160.075 ;
    END
  END wd_in[496]
  PIN wd_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.705 0.070 1160.775 ;
    END
  END wd_in[497]
  PIN wd_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1161.405 0.070 1161.475 ;
    END
  END wd_in[498]
  PIN wd_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.105 0.070 1162.175 ;
    END
  END wd_in[499]
  PIN wd_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.805 0.070 1162.875 ;
    END
  END wd_in[500]
  PIN wd_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1163.505 0.070 1163.575 ;
    END
  END wd_in[501]
  PIN wd_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.205 0.070 1164.275 ;
    END
  END wd_in[502]
  PIN wd_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.905 0.070 1164.975 ;
    END
  END wd_in[503]
  PIN wd_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.605 0.070 1165.675 ;
    END
  END wd_in[504]
  PIN wd_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1166.305 0.070 1166.375 ;
    END
  END wd_in[505]
  PIN wd_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.005 0.070 1167.075 ;
    END
  END wd_in[506]
  PIN wd_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.705 0.070 1167.775 ;
    END
  END wd_in[507]
  PIN wd_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1168.405 0.070 1168.475 ;
    END
  END wd_in[508]
  PIN wd_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.105 0.070 1169.175 ;
    END
  END wd_in[509]
  PIN wd_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.805 0.070 1169.875 ;
    END
  END wd_in[510]
  PIN wd_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1170.505 0.070 1170.575 ;
    END
  END wd_in[511]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.525 0.070 1218.595 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.225 0.070 1219.295 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.925 0.070 1219.995 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1220.625 0.070 1220.695 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1221.325 0.070 1221.395 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.025 0.070 1222.095 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.725 0.070 1222.795 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.425 0.070 1223.495 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.125 0.070 1224.195 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.825 0.070 1224.895 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1225.525 0.070 1225.595 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1226.225 0.070 1226.295 ;
    END
  END addr_in[11]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.245 0.070 1274.315 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.945 0.070 1275.015 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1275.645 0.070 1275.715 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 1279.600 ;
      RECT 3.500 1.400 3.780 1279.600 ;
      RECT 5.740 1.400 6.020 1279.600 ;
      RECT 7.980 1.400 8.260 1279.600 ;
      RECT 10.220 1.400 10.500 1279.600 ;
      RECT 12.460 1.400 12.740 1279.600 ;
      RECT 14.700 1.400 14.980 1279.600 ;
      RECT 16.940 1.400 17.220 1279.600 ;
      RECT 19.180 1.400 19.460 1279.600 ;
      RECT 21.420 1.400 21.700 1279.600 ;
      RECT 23.660 1.400 23.940 1279.600 ;
      RECT 25.900 1.400 26.180 1279.600 ;
      RECT 28.140 1.400 28.420 1279.600 ;
      RECT 30.380 1.400 30.660 1279.600 ;
      RECT 32.620 1.400 32.900 1279.600 ;
      RECT 34.860 1.400 35.140 1279.600 ;
      RECT 37.100 1.400 37.380 1279.600 ;
      RECT 39.340 1.400 39.620 1279.600 ;
      RECT 41.580 1.400 41.860 1279.600 ;
      RECT 43.820 1.400 44.100 1279.600 ;
      RECT 46.060 1.400 46.340 1279.600 ;
      RECT 48.300 1.400 48.580 1279.600 ;
      RECT 50.540 1.400 50.820 1279.600 ;
      RECT 52.780 1.400 53.060 1279.600 ;
      RECT 55.020 1.400 55.300 1279.600 ;
      RECT 57.260 1.400 57.540 1279.600 ;
      RECT 59.500 1.400 59.780 1279.600 ;
      RECT 61.740 1.400 62.020 1279.600 ;
      RECT 63.980 1.400 64.260 1279.600 ;
      RECT 66.220 1.400 66.500 1279.600 ;
      RECT 68.460 1.400 68.740 1279.600 ;
      RECT 70.700 1.400 70.980 1279.600 ;
      RECT 72.940 1.400 73.220 1279.600 ;
      RECT 75.180 1.400 75.460 1279.600 ;
      RECT 77.420 1.400 77.700 1279.600 ;
      RECT 79.660 1.400 79.940 1279.600 ;
      RECT 81.900 1.400 82.180 1279.600 ;
      RECT 84.140 1.400 84.420 1279.600 ;
      RECT 86.380 1.400 86.660 1279.600 ;
      RECT 88.620 1.400 88.900 1279.600 ;
      RECT 90.860 1.400 91.140 1279.600 ;
      RECT 93.100 1.400 93.380 1279.600 ;
      RECT 95.340 1.400 95.620 1279.600 ;
      RECT 97.580 1.400 97.860 1279.600 ;
      RECT 99.820 1.400 100.100 1279.600 ;
      RECT 102.060 1.400 102.340 1279.600 ;
      RECT 104.300 1.400 104.580 1279.600 ;
      RECT 106.540 1.400 106.820 1279.600 ;
      RECT 108.780 1.400 109.060 1279.600 ;
      RECT 111.020 1.400 111.300 1279.600 ;
      RECT 113.260 1.400 113.540 1279.600 ;
      RECT 115.500 1.400 115.780 1279.600 ;
      RECT 117.740 1.400 118.020 1279.600 ;
      RECT 119.980 1.400 120.260 1279.600 ;
      RECT 122.220 1.400 122.500 1279.600 ;
      RECT 124.460 1.400 124.740 1279.600 ;
      RECT 126.700 1.400 126.980 1279.600 ;
      RECT 128.940 1.400 129.220 1279.600 ;
      RECT 131.180 1.400 131.460 1279.600 ;
      RECT 133.420 1.400 133.700 1279.600 ;
      RECT 135.660 1.400 135.940 1279.600 ;
      RECT 137.900 1.400 138.180 1279.600 ;
      RECT 140.140 1.400 140.420 1279.600 ;
      RECT 142.380 1.400 142.660 1279.600 ;
      RECT 144.620 1.400 144.900 1279.600 ;
      RECT 146.860 1.400 147.140 1279.600 ;
      RECT 149.100 1.400 149.380 1279.600 ;
      RECT 151.340 1.400 151.620 1279.600 ;
      RECT 153.580 1.400 153.860 1279.600 ;
      RECT 155.820 1.400 156.100 1279.600 ;
      RECT 158.060 1.400 158.340 1279.600 ;
      RECT 160.300 1.400 160.580 1279.600 ;
      RECT 162.540 1.400 162.820 1279.600 ;
      RECT 164.780 1.400 165.060 1279.600 ;
      RECT 167.020 1.400 167.300 1279.600 ;
      RECT 169.260 1.400 169.540 1279.600 ;
      RECT 171.500 1.400 171.780 1279.600 ;
      RECT 173.740 1.400 174.020 1279.600 ;
      RECT 175.980 1.400 176.260 1279.600 ;
      RECT 178.220 1.400 178.500 1279.600 ;
      RECT 180.460 1.400 180.740 1279.600 ;
      RECT 182.700 1.400 182.980 1279.600 ;
      RECT 184.940 1.400 185.220 1279.600 ;
      RECT 187.180 1.400 187.460 1279.600 ;
      RECT 189.420 1.400 189.700 1279.600 ;
      RECT 191.660 1.400 191.940 1279.600 ;
      RECT 193.900 1.400 194.180 1279.600 ;
      RECT 196.140 1.400 196.420 1279.600 ;
      RECT 198.380 1.400 198.660 1279.600 ;
      RECT 200.620 1.400 200.900 1279.600 ;
      RECT 202.860 1.400 203.140 1279.600 ;
      RECT 205.100 1.400 205.380 1279.600 ;
      RECT 207.340 1.400 207.620 1279.600 ;
      RECT 209.580 1.400 209.860 1279.600 ;
      RECT 211.820 1.400 212.100 1279.600 ;
      RECT 214.060 1.400 214.340 1279.600 ;
      RECT 216.300 1.400 216.580 1279.600 ;
      RECT 218.540 1.400 218.820 1279.600 ;
      RECT 220.780 1.400 221.060 1279.600 ;
      RECT 223.020 1.400 223.300 1279.600 ;
      RECT 225.260 1.400 225.540 1279.600 ;
      RECT 227.500 1.400 227.780 1279.600 ;
      RECT 229.740 1.400 230.020 1279.600 ;
      RECT 231.980 1.400 232.260 1279.600 ;
      RECT 234.220 1.400 234.500 1279.600 ;
      RECT 236.460 1.400 236.740 1279.600 ;
      RECT 238.700 1.400 238.980 1279.600 ;
      RECT 240.940 1.400 241.220 1279.600 ;
      RECT 243.180 1.400 243.460 1279.600 ;
      RECT 245.420 1.400 245.700 1279.600 ;
      RECT 247.660 1.400 247.940 1279.600 ;
      RECT 249.900 1.400 250.180 1279.600 ;
      RECT 252.140 1.400 252.420 1279.600 ;
      RECT 254.380 1.400 254.660 1279.600 ;
      RECT 256.620 1.400 256.900 1279.600 ;
      RECT 258.860 1.400 259.140 1279.600 ;
      RECT 261.100 1.400 261.380 1279.600 ;
      RECT 263.340 1.400 263.620 1279.600 ;
      RECT 265.580 1.400 265.860 1279.600 ;
      RECT 267.820 1.400 268.100 1279.600 ;
      RECT 270.060 1.400 270.340 1279.600 ;
      RECT 272.300 1.400 272.580 1279.600 ;
      RECT 274.540 1.400 274.820 1279.600 ;
      RECT 276.780 1.400 277.060 1279.600 ;
      RECT 279.020 1.400 279.300 1279.600 ;
      RECT 281.260 1.400 281.540 1279.600 ;
      RECT 283.500 1.400 283.780 1279.600 ;
      RECT 285.740 1.400 286.020 1279.600 ;
      RECT 287.980 1.400 288.260 1279.600 ;
      RECT 290.220 1.400 290.500 1279.600 ;
      RECT 292.460 1.400 292.740 1279.600 ;
      RECT 294.700 1.400 294.980 1279.600 ;
      RECT 296.940 1.400 297.220 1279.600 ;
      RECT 299.180 1.400 299.460 1279.600 ;
      RECT 301.420 1.400 301.700 1279.600 ;
      RECT 303.660 1.400 303.940 1279.600 ;
      RECT 305.900 1.400 306.180 1279.600 ;
      RECT 308.140 1.400 308.420 1279.600 ;
      RECT 310.380 1.400 310.660 1279.600 ;
      RECT 312.620 1.400 312.900 1279.600 ;
      RECT 314.860 1.400 315.140 1279.600 ;
      RECT 317.100 1.400 317.380 1279.600 ;
      RECT 319.340 1.400 319.620 1279.600 ;
      RECT 321.580 1.400 321.860 1279.600 ;
      RECT 323.820 1.400 324.100 1279.600 ;
      RECT 326.060 1.400 326.340 1279.600 ;
      RECT 328.300 1.400 328.580 1279.600 ;
      RECT 330.540 1.400 330.820 1279.600 ;
      RECT 332.780 1.400 333.060 1279.600 ;
      RECT 335.020 1.400 335.300 1279.600 ;
      RECT 337.260 1.400 337.540 1279.600 ;
      RECT 339.500 1.400 339.780 1279.600 ;
      RECT 341.740 1.400 342.020 1279.600 ;
      RECT 343.980 1.400 344.260 1279.600 ;
      RECT 346.220 1.400 346.500 1279.600 ;
      RECT 348.460 1.400 348.740 1279.600 ;
      RECT 350.700 1.400 350.980 1279.600 ;
      RECT 352.940 1.400 353.220 1279.600 ;
      RECT 355.180 1.400 355.460 1279.600 ;
      RECT 357.420 1.400 357.700 1279.600 ;
      RECT 359.660 1.400 359.940 1279.600 ;
      RECT 361.900 1.400 362.180 1279.600 ;
      RECT 364.140 1.400 364.420 1279.600 ;
      RECT 366.380 1.400 366.660 1279.600 ;
      RECT 368.620 1.400 368.900 1279.600 ;
      RECT 370.860 1.400 371.140 1279.600 ;
      RECT 373.100 1.400 373.380 1279.600 ;
      RECT 375.340 1.400 375.620 1279.600 ;
      RECT 377.580 1.400 377.860 1279.600 ;
      RECT 379.820 1.400 380.100 1279.600 ;
      RECT 382.060 1.400 382.340 1279.600 ;
      RECT 384.300 1.400 384.580 1279.600 ;
      RECT 386.540 1.400 386.820 1279.600 ;
      RECT 388.780 1.400 389.060 1279.600 ;
      RECT 391.020 1.400 391.300 1279.600 ;
      RECT 393.260 1.400 393.540 1279.600 ;
      RECT 395.500 1.400 395.780 1279.600 ;
      RECT 397.740 1.400 398.020 1279.600 ;
      RECT 399.980 1.400 400.260 1279.600 ;
      RECT 402.220 1.400 402.500 1279.600 ;
      RECT 404.460 1.400 404.740 1279.600 ;
      RECT 406.700 1.400 406.980 1279.600 ;
      RECT 408.940 1.400 409.220 1279.600 ;
      RECT 411.180 1.400 411.460 1279.600 ;
      RECT 413.420 1.400 413.700 1279.600 ;
      RECT 415.660 1.400 415.940 1279.600 ;
      RECT 417.900 1.400 418.180 1279.600 ;
      RECT 420.140 1.400 420.420 1279.600 ;
      RECT 422.380 1.400 422.660 1279.600 ;
      RECT 424.620 1.400 424.900 1279.600 ;
      RECT 426.860 1.400 427.140 1279.600 ;
      RECT 429.100 1.400 429.380 1279.600 ;
      RECT 431.340 1.400 431.620 1279.600 ;
      RECT 433.580 1.400 433.860 1279.600 ;
      RECT 435.820 1.400 436.100 1279.600 ;
      RECT 438.060 1.400 438.340 1279.600 ;
      RECT 440.300 1.400 440.580 1279.600 ;
      RECT 442.540 1.400 442.820 1279.600 ;
      RECT 444.780 1.400 445.060 1279.600 ;
      RECT 447.020 1.400 447.300 1279.600 ;
      RECT 449.260 1.400 449.540 1279.600 ;
      RECT 451.500 1.400 451.780 1279.600 ;
      RECT 453.740 1.400 454.020 1279.600 ;
      RECT 455.980 1.400 456.260 1279.600 ;
      RECT 458.220 1.400 458.500 1279.600 ;
      RECT 460.460 1.400 460.740 1279.600 ;
      RECT 462.700 1.400 462.980 1279.600 ;
      RECT 464.940 1.400 465.220 1279.600 ;
      RECT 467.180 1.400 467.460 1279.600 ;
      RECT 469.420 1.400 469.700 1279.600 ;
      RECT 471.660 1.400 471.940 1279.600 ;
      RECT 473.900 1.400 474.180 1279.600 ;
      RECT 476.140 1.400 476.420 1279.600 ;
      RECT 478.380 1.400 478.660 1279.600 ;
      RECT 480.620 1.400 480.900 1279.600 ;
      RECT 482.860 1.400 483.140 1279.600 ;
      RECT 485.100 1.400 485.380 1279.600 ;
      RECT 487.340 1.400 487.620 1279.600 ;
      RECT 489.580 1.400 489.860 1279.600 ;
      RECT 491.820 1.400 492.100 1279.600 ;
      RECT 494.060 1.400 494.340 1279.600 ;
      RECT 496.300 1.400 496.580 1279.600 ;
      RECT 498.540 1.400 498.820 1279.600 ;
      RECT 500.780 1.400 501.060 1279.600 ;
      RECT 503.020 1.400 503.300 1279.600 ;
      RECT 505.260 1.400 505.540 1279.600 ;
      RECT 507.500 1.400 507.780 1279.600 ;
      RECT 509.740 1.400 510.020 1279.600 ;
      RECT 511.980 1.400 512.260 1279.600 ;
      RECT 514.220 1.400 514.500 1279.600 ;
      RECT 516.460 1.400 516.740 1279.600 ;
      RECT 518.700 1.400 518.980 1279.600 ;
      RECT 520.940 1.400 521.220 1279.600 ;
      RECT 523.180 1.400 523.460 1279.600 ;
      RECT 525.420 1.400 525.700 1279.600 ;
      RECT 527.660 1.400 527.940 1279.600 ;
      RECT 529.900 1.400 530.180 1279.600 ;
      RECT 532.140 1.400 532.420 1279.600 ;
      RECT 534.380 1.400 534.660 1279.600 ;
      RECT 536.620 1.400 536.900 1279.600 ;
      RECT 538.860 1.400 539.140 1279.600 ;
      RECT 541.100 1.400 541.380 1279.600 ;
      RECT 543.340 1.400 543.620 1279.600 ;
      RECT 545.580 1.400 545.860 1279.600 ;
      RECT 547.820 1.400 548.100 1279.600 ;
      RECT 550.060 1.400 550.340 1279.600 ;
      RECT 552.300 1.400 552.580 1279.600 ;
      RECT 554.540 1.400 554.820 1279.600 ;
      RECT 556.780 1.400 557.060 1279.600 ;
      RECT 559.020 1.400 559.300 1279.600 ;
      RECT 561.260 1.400 561.540 1279.600 ;
      RECT 563.500 1.400 563.780 1279.600 ;
      RECT 565.740 1.400 566.020 1279.600 ;
      RECT 567.980 1.400 568.260 1279.600 ;
      RECT 570.220 1.400 570.500 1279.600 ;
      RECT 572.460 1.400 572.740 1279.600 ;
      RECT 574.700 1.400 574.980 1279.600 ;
      RECT 576.940 1.400 577.220 1279.600 ;
      RECT 579.180 1.400 579.460 1279.600 ;
      RECT 581.420 1.400 581.700 1279.600 ;
      RECT 583.660 1.400 583.940 1279.600 ;
      RECT 585.900 1.400 586.180 1279.600 ;
      RECT 588.140 1.400 588.420 1279.600 ;
      RECT 590.380 1.400 590.660 1279.600 ;
      RECT 592.620 1.400 592.900 1279.600 ;
      RECT 594.860 1.400 595.140 1279.600 ;
      RECT 597.100 1.400 597.380 1279.600 ;
      RECT 599.340 1.400 599.620 1279.600 ;
      RECT 601.580 1.400 601.860 1279.600 ;
      RECT 603.820 1.400 604.100 1279.600 ;
      RECT 606.060 1.400 606.340 1279.600 ;
      RECT 608.300 1.400 608.580 1279.600 ;
      RECT 610.540 1.400 610.820 1279.600 ;
      RECT 612.780 1.400 613.060 1279.600 ;
      RECT 615.020 1.400 615.300 1279.600 ;
      RECT 617.260 1.400 617.540 1279.600 ;
      RECT 619.500 1.400 619.780 1279.600 ;
      RECT 621.740 1.400 622.020 1279.600 ;
      RECT 623.980 1.400 624.260 1279.600 ;
      RECT 626.220 1.400 626.500 1279.600 ;
      RECT 628.460 1.400 628.740 1279.600 ;
      RECT 630.700 1.400 630.980 1279.600 ;
      RECT 632.940 1.400 633.220 1279.600 ;
      RECT 635.180 1.400 635.460 1279.600 ;
      RECT 637.420 1.400 637.700 1279.600 ;
      RECT 639.660 1.400 639.940 1279.600 ;
      RECT 641.900 1.400 642.180 1279.600 ;
      RECT 644.140 1.400 644.420 1279.600 ;
      RECT 646.380 1.400 646.660 1279.600 ;
      RECT 648.620 1.400 648.900 1279.600 ;
      RECT 650.860 1.400 651.140 1279.600 ;
      RECT 653.100 1.400 653.380 1279.600 ;
      RECT 655.340 1.400 655.620 1279.600 ;
      RECT 657.580 1.400 657.860 1279.600 ;
      RECT 659.820 1.400 660.100 1279.600 ;
      RECT 662.060 1.400 662.340 1279.600 ;
      RECT 664.300 1.400 664.580 1279.600 ;
      RECT 666.540 1.400 666.820 1279.600 ;
      RECT 668.780 1.400 669.060 1279.600 ;
      RECT 671.020 1.400 671.300 1279.600 ;
      RECT 673.260 1.400 673.540 1279.600 ;
      RECT 675.500 1.400 675.780 1279.600 ;
      RECT 677.740 1.400 678.020 1279.600 ;
      RECT 679.980 1.400 680.260 1279.600 ;
      RECT 682.220 1.400 682.500 1279.600 ;
      RECT 684.460 1.400 684.740 1279.600 ;
      RECT 686.700 1.400 686.980 1279.600 ;
      RECT 688.940 1.400 689.220 1279.600 ;
      RECT 691.180 1.400 691.460 1279.600 ;
      RECT 693.420 1.400 693.700 1279.600 ;
      RECT 695.660 1.400 695.940 1279.600 ;
      RECT 697.900 1.400 698.180 1279.600 ;
      RECT 700.140 1.400 700.420 1279.600 ;
      RECT 702.380 1.400 702.660 1279.600 ;
      RECT 704.620 1.400 704.900 1279.600 ;
      RECT 706.860 1.400 707.140 1279.600 ;
      RECT 709.100 1.400 709.380 1279.600 ;
      RECT 711.340 1.400 711.620 1279.600 ;
      RECT 713.580 1.400 713.860 1279.600 ;
      RECT 715.820 1.400 716.100 1279.600 ;
      RECT 718.060 1.400 718.340 1279.600 ;
      RECT 720.300 1.400 720.580 1279.600 ;
      RECT 722.540 1.400 722.820 1279.600 ;
      RECT 724.780 1.400 725.060 1279.600 ;
      RECT 727.020 1.400 727.300 1279.600 ;
      RECT 729.260 1.400 729.540 1279.600 ;
      RECT 731.500 1.400 731.780 1279.600 ;
      RECT 733.740 1.400 734.020 1279.600 ;
      RECT 735.980 1.400 736.260 1279.600 ;
      RECT 738.220 1.400 738.500 1279.600 ;
      RECT 740.460 1.400 740.740 1279.600 ;
      RECT 742.700 1.400 742.980 1279.600 ;
      RECT 744.940 1.400 745.220 1279.600 ;
      RECT 747.180 1.400 747.460 1279.600 ;
      RECT 749.420 1.400 749.700 1279.600 ;
      RECT 751.660 1.400 751.940 1279.600 ;
      RECT 753.900 1.400 754.180 1279.600 ;
      RECT 756.140 1.400 756.420 1279.600 ;
      RECT 758.380 1.400 758.660 1279.600 ;
      RECT 760.620 1.400 760.900 1279.600 ;
      RECT 762.860 1.400 763.140 1279.600 ;
      RECT 765.100 1.400 765.380 1279.600 ;
      RECT 767.340 1.400 767.620 1279.600 ;
      RECT 769.580 1.400 769.860 1279.600 ;
      RECT 771.820 1.400 772.100 1279.600 ;
      RECT 774.060 1.400 774.340 1279.600 ;
      RECT 776.300 1.400 776.580 1279.600 ;
      RECT 778.540 1.400 778.820 1279.600 ;
      RECT 780.780 1.400 781.060 1279.600 ;
      RECT 783.020 1.400 783.300 1279.600 ;
      RECT 785.260 1.400 785.540 1279.600 ;
      RECT 787.500 1.400 787.780 1279.600 ;
      RECT 789.740 1.400 790.020 1279.600 ;
      RECT 791.980 1.400 792.260 1279.600 ;
      RECT 794.220 1.400 794.500 1279.600 ;
      RECT 796.460 1.400 796.740 1279.600 ;
      RECT 798.700 1.400 798.980 1279.600 ;
      RECT 800.940 1.400 801.220 1279.600 ;
      RECT 803.180 1.400 803.460 1279.600 ;
      RECT 805.420 1.400 805.700 1279.600 ;
      RECT 807.660 1.400 807.940 1279.600 ;
      RECT 809.900 1.400 810.180 1279.600 ;
      RECT 812.140 1.400 812.420 1279.600 ;
      RECT 814.380 1.400 814.660 1279.600 ;
      RECT 816.620 1.400 816.900 1279.600 ;
      RECT 818.860 1.400 819.140 1279.600 ;
      RECT 821.100 1.400 821.380 1279.600 ;
      RECT 823.340 1.400 823.620 1279.600 ;
      RECT 825.580 1.400 825.860 1279.600 ;
      RECT 827.820 1.400 828.100 1279.600 ;
      RECT 830.060 1.400 830.340 1279.600 ;
      RECT 832.300 1.400 832.580 1279.600 ;
      RECT 834.540 1.400 834.820 1279.600 ;
      RECT 836.780 1.400 837.060 1279.600 ;
      RECT 839.020 1.400 839.300 1279.600 ;
      RECT 841.260 1.400 841.540 1279.600 ;
      RECT 843.500 1.400 843.780 1279.600 ;
      RECT 845.740 1.400 846.020 1279.600 ;
      RECT 847.980 1.400 848.260 1279.600 ;
      RECT 850.220 1.400 850.500 1279.600 ;
      RECT 852.460 1.400 852.740 1279.600 ;
      RECT 854.700 1.400 854.980 1279.600 ;
      RECT 856.940 1.400 857.220 1279.600 ;
      RECT 859.180 1.400 859.460 1279.600 ;
      RECT 861.420 1.400 861.700 1279.600 ;
      RECT 863.660 1.400 863.940 1279.600 ;
      RECT 865.900 1.400 866.180 1279.600 ;
      RECT 868.140 1.400 868.420 1279.600 ;
      RECT 870.380 1.400 870.660 1279.600 ;
      RECT 872.620 1.400 872.900 1279.600 ;
      RECT 874.860 1.400 875.140 1279.600 ;
      RECT 877.100 1.400 877.380 1279.600 ;
      RECT 879.340 1.400 879.620 1279.600 ;
      RECT 881.580 1.400 881.860 1279.600 ;
      RECT 883.820 1.400 884.100 1279.600 ;
      RECT 886.060 1.400 886.340 1279.600 ;
      RECT 888.300 1.400 888.580 1279.600 ;
      RECT 890.540 1.400 890.820 1279.600 ;
      RECT 892.780 1.400 893.060 1279.600 ;
      RECT 895.020 1.400 895.300 1279.600 ;
      RECT 897.260 1.400 897.540 1279.600 ;
      RECT 899.500 1.400 899.780 1279.600 ;
      RECT 901.740 1.400 902.020 1279.600 ;
      RECT 903.980 1.400 904.260 1279.600 ;
      RECT 906.220 1.400 906.500 1279.600 ;
      RECT 908.460 1.400 908.740 1279.600 ;
      RECT 910.700 1.400 910.980 1279.600 ;
      RECT 912.940 1.400 913.220 1279.600 ;
      RECT 915.180 1.400 915.460 1279.600 ;
      RECT 917.420 1.400 917.700 1279.600 ;
      RECT 919.660 1.400 919.940 1279.600 ;
      RECT 921.900 1.400 922.180 1279.600 ;
      RECT 924.140 1.400 924.420 1279.600 ;
      RECT 926.380 1.400 926.660 1279.600 ;
      RECT 928.620 1.400 928.900 1279.600 ;
      RECT 930.860 1.400 931.140 1279.600 ;
      RECT 933.100 1.400 933.380 1279.600 ;
      RECT 935.340 1.400 935.620 1279.600 ;
      RECT 937.580 1.400 937.860 1279.600 ;
      RECT 939.820 1.400 940.100 1279.600 ;
      RECT 942.060 1.400 942.340 1279.600 ;
      RECT 944.300 1.400 944.580 1279.600 ;
      RECT 946.540 1.400 946.820 1279.600 ;
      RECT 948.780 1.400 949.060 1279.600 ;
      RECT 951.020 1.400 951.300 1279.600 ;
      RECT 953.260 1.400 953.540 1279.600 ;
      RECT 955.500 1.400 955.780 1279.600 ;
      RECT 957.740 1.400 958.020 1279.600 ;
      RECT 959.980 1.400 960.260 1279.600 ;
      RECT 962.220 1.400 962.500 1279.600 ;
      RECT 964.460 1.400 964.740 1279.600 ;
      RECT 966.700 1.400 966.980 1279.600 ;
      RECT 968.940 1.400 969.220 1279.600 ;
      RECT 971.180 1.400 971.460 1279.600 ;
      RECT 973.420 1.400 973.700 1279.600 ;
      RECT 975.660 1.400 975.940 1279.600 ;
      RECT 977.900 1.400 978.180 1279.600 ;
      RECT 980.140 1.400 980.420 1279.600 ;
      RECT 982.380 1.400 982.660 1279.600 ;
      RECT 984.620 1.400 984.900 1279.600 ;
      RECT 986.860 1.400 987.140 1279.600 ;
      RECT 989.100 1.400 989.380 1279.600 ;
      RECT 991.340 1.400 991.620 1279.600 ;
      RECT 993.580 1.400 993.860 1279.600 ;
      RECT 995.820 1.400 996.100 1279.600 ;
      RECT 998.060 1.400 998.340 1279.600 ;
      RECT 1000.300 1.400 1000.580 1279.600 ;
      RECT 1002.540 1.400 1002.820 1279.600 ;
      RECT 1004.780 1.400 1005.060 1279.600 ;
      RECT 1007.020 1.400 1007.300 1279.600 ;
      RECT 1009.260 1.400 1009.540 1279.600 ;
      RECT 1011.500 1.400 1011.780 1279.600 ;
      RECT 1013.740 1.400 1014.020 1279.600 ;
      RECT 1015.980 1.400 1016.260 1279.600 ;
      RECT 1018.220 1.400 1018.500 1279.600 ;
      RECT 1020.460 1.400 1020.740 1279.600 ;
      RECT 1022.700 1.400 1022.980 1279.600 ;
      RECT 1024.940 1.400 1025.220 1279.600 ;
      RECT 1027.180 1.400 1027.460 1279.600 ;
      RECT 1029.420 1.400 1029.700 1279.600 ;
      RECT 1031.660 1.400 1031.940 1279.600 ;
      RECT 1033.900 1.400 1034.180 1279.600 ;
      RECT 1036.140 1.400 1036.420 1279.600 ;
      RECT 1038.380 1.400 1038.660 1279.600 ;
      RECT 1040.620 1.400 1040.900 1279.600 ;
      RECT 1042.860 1.400 1043.140 1279.600 ;
      RECT 1045.100 1.400 1045.380 1279.600 ;
      RECT 1047.340 1.400 1047.620 1279.600 ;
      RECT 1049.580 1.400 1049.860 1279.600 ;
      RECT 1051.820 1.400 1052.100 1279.600 ;
      RECT 1054.060 1.400 1054.340 1279.600 ;
      RECT 1056.300 1.400 1056.580 1279.600 ;
      RECT 1058.540 1.400 1058.820 1279.600 ;
      RECT 1060.780 1.400 1061.060 1279.600 ;
      RECT 1063.020 1.400 1063.300 1279.600 ;
      RECT 1065.260 1.400 1065.540 1279.600 ;
      RECT 1067.500 1.400 1067.780 1279.600 ;
      RECT 1069.740 1.400 1070.020 1279.600 ;
      RECT 1071.980 1.400 1072.260 1279.600 ;
      RECT 1074.220 1.400 1074.500 1279.600 ;
      RECT 1076.460 1.400 1076.740 1279.600 ;
      RECT 1078.700 1.400 1078.980 1279.600 ;
      RECT 1080.940 1.400 1081.220 1279.600 ;
      RECT 1083.180 1.400 1083.460 1279.600 ;
      RECT 1085.420 1.400 1085.700 1279.600 ;
      RECT 1087.660 1.400 1087.940 1279.600 ;
      RECT 1089.900 1.400 1090.180 1279.600 ;
      RECT 1092.140 1.400 1092.420 1279.600 ;
      RECT 1094.380 1.400 1094.660 1279.600 ;
      RECT 1096.620 1.400 1096.900 1279.600 ;
      RECT 1098.860 1.400 1099.140 1279.600 ;
      RECT 1101.100 1.400 1101.380 1279.600 ;
      RECT 1103.340 1.400 1103.620 1279.600 ;
      RECT 1105.580 1.400 1105.860 1279.600 ;
      RECT 1107.820 1.400 1108.100 1279.600 ;
      RECT 1110.060 1.400 1110.340 1279.600 ;
      RECT 1112.300 1.400 1112.580 1279.600 ;
      RECT 1114.540 1.400 1114.820 1279.600 ;
      RECT 1116.780 1.400 1117.060 1279.600 ;
      RECT 1119.020 1.400 1119.300 1279.600 ;
      RECT 1121.260 1.400 1121.540 1279.600 ;
      RECT 1123.500 1.400 1123.780 1279.600 ;
      RECT 1125.740 1.400 1126.020 1279.600 ;
      RECT 1127.980 1.400 1128.260 1279.600 ;
      RECT 1130.220 1.400 1130.500 1279.600 ;
      RECT 1132.460 1.400 1132.740 1279.600 ;
      RECT 1134.700 1.400 1134.980 1279.600 ;
      RECT 1136.940 1.400 1137.220 1279.600 ;
      RECT 1139.180 1.400 1139.460 1279.600 ;
      RECT 1141.420 1.400 1141.700 1279.600 ;
      RECT 1143.660 1.400 1143.940 1279.600 ;
      RECT 1145.900 1.400 1146.180 1279.600 ;
      RECT 1148.140 1.400 1148.420 1279.600 ;
      RECT 1150.380 1.400 1150.660 1279.600 ;
      RECT 1152.620 1.400 1152.900 1279.600 ;
      RECT 1154.860 1.400 1155.140 1279.600 ;
      RECT 1157.100 1.400 1157.380 1279.600 ;
      RECT 1159.340 1.400 1159.620 1279.600 ;
      RECT 1161.580 1.400 1161.860 1279.600 ;
      RECT 1163.820 1.400 1164.100 1279.600 ;
      RECT 1166.060 1.400 1166.340 1279.600 ;
      RECT 1168.300 1.400 1168.580 1279.600 ;
      RECT 1170.540 1.400 1170.820 1279.600 ;
      RECT 1172.780 1.400 1173.060 1279.600 ;
      RECT 1175.020 1.400 1175.300 1279.600 ;
      RECT 1177.260 1.400 1177.540 1279.600 ;
      RECT 1179.500 1.400 1179.780 1279.600 ;
      RECT 1181.740 1.400 1182.020 1279.600 ;
      RECT 1183.980 1.400 1184.260 1279.600 ;
      RECT 1186.220 1.400 1186.500 1279.600 ;
      RECT 1188.460 1.400 1188.740 1279.600 ;
      RECT 1190.700 1.400 1190.980 1279.600 ;
      RECT 1192.940 1.400 1193.220 1279.600 ;
      RECT 1195.180 1.400 1195.460 1279.600 ;
      RECT 1197.420 1.400 1197.700 1279.600 ;
      RECT 1199.660 1.400 1199.940 1279.600 ;
      RECT 1201.900 1.400 1202.180 1279.600 ;
      RECT 1204.140 1.400 1204.420 1279.600 ;
      RECT 1206.380 1.400 1206.660 1279.600 ;
      RECT 1208.620 1.400 1208.900 1279.600 ;
      RECT 1210.860 1.400 1211.140 1279.600 ;
      RECT 1213.100 1.400 1213.380 1279.600 ;
      RECT 1215.340 1.400 1215.620 1279.600 ;
      RECT 1217.580 1.400 1217.860 1279.600 ;
      RECT 1219.820 1.400 1220.100 1279.600 ;
      RECT 1222.060 1.400 1222.340 1279.600 ;
      RECT 1224.300 1.400 1224.580 1279.600 ;
      RECT 1226.540 1.400 1226.820 1279.600 ;
      RECT 1228.780 1.400 1229.060 1279.600 ;
      RECT 1231.020 1.400 1231.300 1279.600 ;
      RECT 1233.260 1.400 1233.540 1279.600 ;
      RECT 1235.500 1.400 1235.780 1279.600 ;
      RECT 1237.740 1.400 1238.020 1279.600 ;
      RECT 1239.980 1.400 1240.260 1279.600 ;
      RECT 1242.220 1.400 1242.500 1279.600 ;
      RECT 1244.460 1.400 1244.740 1279.600 ;
      RECT 1246.700 1.400 1246.980 1279.600 ;
      RECT 1248.940 1.400 1249.220 1279.600 ;
      RECT 1251.180 1.400 1251.460 1279.600 ;
      RECT 1253.420 1.400 1253.700 1279.600 ;
      RECT 1255.660 1.400 1255.940 1279.600 ;
      RECT 1257.900 1.400 1258.180 1279.600 ;
      RECT 1260.140 1.400 1260.420 1279.600 ;
      RECT 1262.380 1.400 1262.660 1279.600 ;
      RECT 1264.620 1.400 1264.900 1279.600 ;
      RECT 1266.860 1.400 1267.140 1279.600 ;
      RECT 1269.100 1.400 1269.380 1279.600 ;
      RECT 1271.340 1.400 1271.620 1279.600 ;
      RECT 1273.580 1.400 1273.860 1279.600 ;
      RECT 1275.820 1.400 1276.100 1279.600 ;
      RECT 1278.060 1.400 1278.340 1279.600 ;
      RECT 1280.300 1.400 1280.580 1279.600 ;
      RECT 1282.540 1.400 1282.820 1279.600 ;
      RECT 1284.780 1.400 1285.060 1279.600 ;
      RECT 1287.020 1.400 1287.300 1279.600 ;
      RECT 1289.260 1.400 1289.540 1279.600 ;
      RECT 1291.500 1.400 1291.780 1279.600 ;
      RECT 1293.740 1.400 1294.020 1279.600 ;
      RECT 1295.980 1.400 1296.260 1279.600 ;
      RECT 1298.220 1.400 1298.500 1279.600 ;
      RECT 1300.460 1.400 1300.740 1279.600 ;
      RECT 1302.700 1.400 1302.980 1279.600 ;
      RECT 1304.940 1.400 1305.220 1279.600 ;
      RECT 1307.180 1.400 1307.460 1279.600 ;
      RECT 1309.420 1.400 1309.700 1279.600 ;
      RECT 1311.660 1.400 1311.940 1279.600 ;
      RECT 1313.900 1.400 1314.180 1279.600 ;
      RECT 1316.140 1.400 1316.420 1279.600 ;
      RECT 1318.380 1.400 1318.660 1279.600 ;
      RECT 1320.620 1.400 1320.900 1279.600 ;
      RECT 1322.860 1.400 1323.140 1279.600 ;
      RECT 1325.100 1.400 1325.380 1279.600 ;
      RECT 1327.340 1.400 1327.620 1279.600 ;
      RECT 1329.580 1.400 1329.860 1279.600 ;
      RECT 1331.820 1.400 1332.100 1279.600 ;
      RECT 1334.060 1.400 1334.340 1279.600 ;
      RECT 1336.300 1.400 1336.580 1279.600 ;
      RECT 1338.540 1.400 1338.820 1279.600 ;
      RECT 1340.780 1.400 1341.060 1279.600 ;
      RECT 1343.020 1.400 1343.300 1279.600 ;
      RECT 1345.260 1.400 1345.540 1279.600 ;
      RECT 1347.500 1.400 1347.780 1279.600 ;
      RECT 1349.740 1.400 1350.020 1279.600 ;
      RECT 1351.980 1.400 1352.260 1279.600 ;
      RECT 1354.220 1.400 1354.500 1279.600 ;
      RECT 1356.460 1.400 1356.740 1279.600 ;
      RECT 1358.700 1.400 1358.980 1279.600 ;
      RECT 1360.940 1.400 1361.220 1279.600 ;
      RECT 1363.180 1.400 1363.460 1279.600 ;
      RECT 1365.420 1.400 1365.700 1279.600 ;
      RECT 1367.660 1.400 1367.940 1279.600 ;
      RECT 1369.900 1.400 1370.180 1279.600 ;
      RECT 1372.140 1.400 1372.420 1279.600 ;
      RECT 1374.380 1.400 1374.660 1279.600 ;
      RECT 1376.620 1.400 1376.900 1279.600 ;
      RECT 1378.860 1.400 1379.140 1279.600 ;
      RECT 1381.100 1.400 1381.380 1279.600 ;
      RECT 1383.340 1.400 1383.620 1279.600 ;
      RECT 1385.580 1.400 1385.860 1279.600 ;
      RECT 1387.820 1.400 1388.100 1279.600 ;
      RECT 1390.060 1.400 1390.340 1279.600 ;
      RECT 1392.300 1.400 1392.580 1279.600 ;
      RECT 1394.540 1.400 1394.820 1279.600 ;
      RECT 1396.780 1.400 1397.060 1279.600 ;
      RECT 1399.020 1.400 1399.300 1279.600 ;
      RECT 1401.260 1.400 1401.540 1279.600 ;
      RECT 1403.500 1.400 1403.780 1279.600 ;
      RECT 1405.740 1.400 1406.020 1279.600 ;
      RECT 1407.980 1.400 1408.260 1279.600 ;
      RECT 1410.220 1.400 1410.500 1279.600 ;
      RECT 1412.460 1.400 1412.740 1279.600 ;
      RECT 1414.700 1.400 1414.980 1279.600 ;
      RECT 1416.940 1.400 1417.220 1279.600 ;
      RECT 1419.180 1.400 1419.460 1279.600 ;
      RECT 1421.420 1.400 1421.700 1279.600 ;
      RECT 1423.660 1.400 1423.940 1279.600 ;
      RECT 1425.900 1.400 1426.180 1279.600 ;
      RECT 1428.140 1.400 1428.420 1279.600 ;
      RECT 1430.380 1.400 1430.660 1279.600 ;
      RECT 1432.620 1.400 1432.900 1279.600 ;
      RECT 1434.860 1.400 1435.140 1279.600 ;
      RECT 1437.100 1.400 1437.380 1279.600 ;
      RECT 1439.340 1.400 1439.620 1279.600 ;
      RECT 1441.580 1.400 1441.860 1279.600 ;
      RECT 1443.820 1.400 1444.100 1279.600 ;
      RECT 1446.060 1.400 1446.340 1279.600 ;
      RECT 1448.300 1.400 1448.580 1279.600 ;
      RECT 1450.540 1.400 1450.820 1279.600 ;
      RECT 1452.780 1.400 1453.060 1279.600 ;
      RECT 1455.020 1.400 1455.300 1279.600 ;
      RECT 1457.260 1.400 1457.540 1279.600 ;
      RECT 1459.500 1.400 1459.780 1279.600 ;
      RECT 1461.740 1.400 1462.020 1279.600 ;
      RECT 1463.980 1.400 1464.260 1279.600 ;
      RECT 1466.220 1.400 1466.500 1279.600 ;
      RECT 1468.460 1.400 1468.740 1279.600 ;
      RECT 1470.700 1.400 1470.980 1279.600 ;
      RECT 1472.940 1.400 1473.220 1279.600 ;
      RECT 1475.180 1.400 1475.460 1279.600 ;
      RECT 1477.420 1.400 1477.700 1279.600 ;
      RECT 1479.660 1.400 1479.940 1279.600 ;
      RECT 1481.900 1.400 1482.180 1279.600 ;
      RECT 1484.140 1.400 1484.420 1279.600 ;
      RECT 1486.380 1.400 1486.660 1279.600 ;
      RECT 1488.620 1.400 1488.900 1279.600 ;
      RECT 1490.860 1.400 1491.140 1279.600 ;
      RECT 1493.100 1.400 1493.380 1279.600 ;
      RECT 1495.340 1.400 1495.620 1279.600 ;
      RECT 1497.580 1.400 1497.860 1279.600 ;
      RECT 1499.820 1.400 1500.100 1279.600 ;
      RECT 1502.060 1.400 1502.340 1279.600 ;
      RECT 1504.300 1.400 1504.580 1279.600 ;
      RECT 1506.540 1.400 1506.820 1279.600 ;
      RECT 1508.780 1.400 1509.060 1279.600 ;
      RECT 1511.020 1.400 1511.300 1279.600 ;
      RECT 1513.260 1.400 1513.540 1279.600 ;
      RECT 1515.500 1.400 1515.780 1279.600 ;
      RECT 1517.740 1.400 1518.020 1279.600 ;
      RECT 1519.980 1.400 1520.260 1279.600 ;
      RECT 1522.220 1.400 1522.500 1279.600 ;
      RECT 1524.460 1.400 1524.740 1279.600 ;
      RECT 1526.700 1.400 1526.980 1279.600 ;
      RECT 1528.940 1.400 1529.220 1279.600 ;
      RECT 1531.180 1.400 1531.460 1279.600 ;
      RECT 1533.420 1.400 1533.700 1279.600 ;
      RECT 1535.660 1.400 1535.940 1279.600 ;
      RECT 1537.900 1.400 1538.180 1279.600 ;
      RECT 1540.140 1.400 1540.420 1279.600 ;
      RECT 1542.380 1.400 1542.660 1279.600 ;
      RECT 1544.620 1.400 1544.900 1279.600 ;
      RECT 1546.860 1.400 1547.140 1279.600 ;
      RECT 1549.100 1.400 1549.380 1279.600 ;
      RECT 1551.340 1.400 1551.620 1279.600 ;
      RECT 1553.580 1.400 1553.860 1279.600 ;
      RECT 1555.820 1.400 1556.100 1279.600 ;
      RECT 1558.060 1.400 1558.340 1279.600 ;
      RECT 1560.300 1.400 1560.580 1279.600 ;
      RECT 1562.540 1.400 1562.820 1279.600 ;
      RECT 1564.780 1.400 1565.060 1279.600 ;
      RECT 1567.020 1.400 1567.300 1279.600 ;
      RECT 1569.260 1.400 1569.540 1279.600 ;
      RECT 1571.500 1.400 1571.780 1279.600 ;
      RECT 1573.740 1.400 1574.020 1279.600 ;
      RECT 1575.980 1.400 1576.260 1279.600 ;
      RECT 1578.220 1.400 1578.500 1279.600 ;
      RECT 1580.460 1.400 1580.740 1279.600 ;
      RECT 1582.700 1.400 1582.980 1279.600 ;
      RECT 1584.940 1.400 1585.220 1279.600 ;
      RECT 1587.180 1.400 1587.460 1279.600 ;
      RECT 1589.420 1.400 1589.700 1279.600 ;
      RECT 1591.660 1.400 1591.940 1279.600 ;
      RECT 1593.900 1.400 1594.180 1279.600 ;
      RECT 1596.140 1.400 1596.420 1279.600 ;
      RECT 1598.380 1.400 1598.660 1279.600 ;
      RECT 1600.620 1.400 1600.900 1279.600 ;
      RECT 1602.860 1.400 1603.140 1279.600 ;
      RECT 1605.100 1.400 1605.380 1279.600 ;
      RECT 1607.340 1.400 1607.620 1279.600 ;
      RECT 1609.580 1.400 1609.860 1279.600 ;
      RECT 1611.820 1.400 1612.100 1279.600 ;
      RECT 1614.060 1.400 1614.340 1279.600 ;
      RECT 1616.300 1.400 1616.580 1279.600 ;
      RECT 1618.540 1.400 1618.820 1279.600 ;
      RECT 1620.780 1.400 1621.060 1279.600 ;
      RECT 1623.020 1.400 1623.300 1279.600 ;
      RECT 1625.260 1.400 1625.540 1279.600 ;
      RECT 1627.500 1.400 1627.780 1279.600 ;
      RECT 1629.740 1.400 1630.020 1279.600 ;
      RECT 1631.980 1.400 1632.260 1279.600 ;
      RECT 1634.220 1.400 1634.500 1279.600 ;
      RECT 1636.460 1.400 1636.740 1279.600 ;
      RECT 1638.700 1.400 1638.980 1279.600 ;
      RECT 1640.940 1.400 1641.220 1279.600 ;
      RECT 1643.180 1.400 1643.460 1279.600 ;
      RECT 1645.420 1.400 1645.700 1279.600 ;
      RECT 1647.660 1.400 1647.940 1279.600 ;
      RECT 1649.900 1.400 1650.180 1279.600 ;
      RECT 1652.140 1.400 1652.420 1279.600 ;
      RECT 1654.380 1.400 1654.660 1279.600 ;
      RECT 1656.620 1.400 1656.900 1279.600 ;
      RECT 1658.860 1.400 1659.140 1279.600 ;
      RECT 1661.100 1.400 1661.380 1279.600 ;
      RECT 1663.340 1.400 1663.620 1279.600 ;
      RECT 1665.580 1.400 1665.860 1279.600 ;
      RECT 1667.820 1.400 1668.100 1279.600 ;
      RECT 1670.060 1.400 1670.340 1279.600 ;
      RECT 1672.300 1.400 1672.580 1279.600 ;
      RECT 1674.540 1.400 1674.820 1279.600 ;
      RECT 1676.780 1.400 1677.060 1279.600 ;
      RECT 1679.020 1.400 1679.300 1279.600 ;
      RECT 1681.260 1.400 1681.540 1279.600 ;
      RECT 1683.500 1.400 1683.780 1279.600 ;
      RECT 1685.740 1.400 1686.020 1279.600 ;
      RECT 1687.980 1.400 1688.260 1279.600 ;
      RECT 1690.220 1.400 1690.500 1279.600 ;
      RECT 1692.460 1.400 1692.740 1279.600 ;
      RECT 1694.700 1.400 1694.980 1279.600 ;
      RECT 1696.940 1.400 1697.220 1279.600 ;
      RECT 1699.180 1.400 1699.460 1279.600 ;
      RECT 1701.420 1.400 1701.700 1279.600 ;
      RECT 1703.660 1.400 1703.940 1279.600 ;
      RECT 1705.900 1.400 1706.180 1279.600 ;
      RECT 1708.140 1.400 1708.420 1279.600 ;
      RECT 1710.380 1.400 1710.660 1279.600 ;
      RECT 1712.620 1.400 1712.900 1279.600 ;
      RECT 1714.860 1.400 1715.140 1279.600 ;
      RECT 1717.100 1.400 1717.380 1279.600 ;
      RECT 1719.340 1.400 1719.620 1279.600 ;
      RECT 1721.580 1.400 1721.860 1279.600 ;
      RECT 1723.820 1.400 1724.100 1279.600 ;
      RECT 1726.060 1.400 1726.340 1279.600 ;
      RECT 1728.300 1.400 1728.580 1279.600 ;
      RECT 1730.540 1.400 1730.820 1279.600 ;
      RECT 1732.780 1.400 1733.060 1279.600 ;
      RECT 1735.020 1.400 1735.300 1279.600 ;
      RECT 1737.260 1.400 1737.540 1279.600 ;
      RECT 1739.500 1.400 1739.780 1279.600 ;
      RECT 1741.740 1.400 1742.020 1279.600 ;
      RECT 1743.980 1.400 1744.260 1279.600 ;
      RECT 1746.220 1.400 1746.500 1279.600 ;
      RECT 1748.460 1.400 1748.740 1279.600 ;
      RECT 1750.700 1.400 1750.980 1279.600 ;
      RECT 1752.940 1.400 1753.220 1279.600 ;
      RECT 1755.180 1.400 1755.460 1279.600 ;
      RECT 1757.420 1.400 1757.700 1279.600 ;
      RECT 1759.660 1.400 1759.940 1279.600 ;
      RECT 1761.900 1.400 1762.180 1279.600 ;
      RECT 1764.140 1.400 1764.420 1279.600 ;
      RECT 1766.380 1.400 1766.660 1279.600 ;
      RECT 1768.620 1.400 1768.900 1279.600 ;
      RECT 1770.860 1.400 1771.140 1279.600 ;
      RECT 1773.100 1.400 1773.380 1279.600 ;
      RECT 1775.340 1.400 1775.620 1279.600 ;
      RECT 1777.580 1.400 1777.860 1279.600 ;
      RECT 1779.820 1.400 1780.100 1279.600 ;
      RECT 1782.060 1.400 1782.340 1279.600 ;
      RECT 1784.300 1.400 1784.580 1279.600 ;
      RECT 1786.540 1.400 1786.820 1279.600 ;
      RECT 1788.780 1.400 1789.060 1279.600 ;
      RECT 1791.020 1.400 1791.300 1279.600 ;
      RECT 1793.260 1.400 1793.540 1279.600 ;
      RECT 1795.500 1.400 1795.780 1279.600 ;
      RECT 1797.740 1.400 1798.020 1279.600 ;
      RECT 1799.980 1.400 1800.260 1279.600 ;
      RECT 1802.220 1.400 1802.500 1279.600 ;
      RECT 1804.460 1.400 1804.740 1279.600 ;
      RECT 1806.700 1.400 1806.980 1279.600 ;
      RECT 1808.940 1.400 1809.220 1279.600 ;
      RECT 1811.180 1.400 1811.460 1279.600 ;
      RECT 1813.420 1.400 1813.700 1279.600 ;
      RECT 1815.660 1.400 1815.940 1279.600 ;
      RECT 1817.900 1.400 1818.180 1279.600 ;
      RECT 1820.140 1.400 1820.420 1279.600 ;
      RECT 1822.380 1.400 1822.660 1279.600 ;
      RECT 1824.620 1.400 1824.900 1279.600 ;
      RECT 1826.860 1.400 1827.140 1279.600 ;
      RECT 1829.100 1.400 1829.380 1279.600 ;
      RECT 1831.340 1.400 1831.620 1279.600 ;
      RECT 1833.580 1.400 1833.860 1279.600 ;
      RECT 1835.820 1.400 1836.100 1279.600 ;
      RECT 1838.060 1.400 1838.340 1279.600 ;
      RECT 1840.300 1.400 1840.580 1279.600 ;
      RECT 1842.540 1.400 1842.820 1279.600 ;
      RECT 1844.780 1.400 1845.060 1279.600 ;
      RECT 1847.020 1.400 1847.300 1279.600 ;
      RECT 1849.260 1.400 1849.540 1279.600 ;
      RECT 1851.500 1.400 1851.780 1279.600 ;
      RECT 1853.740 1.400 1854.020 1279.600 ;
      RECT 1855.980 1.400 1856.260 1279.600 ;
      RECT 1858.220 1.400 1858.500 1279.600 ;
      RECT 1860.460 1.400 1860.740 1279.600 ;
      RECT 1862.700 1.400 1862.980 1279.600 ;
      RECT 1864.940 1.400 1865.220 1279.600 ;
      RECT 1867.180 1.400 1867.460 1279.600 ;
      RECT 1869.420 1.400 1869.700 1279.600 ;
      RECT 1871.660 1.400 1871.940 1279.600 ;
      RECT 1873.900 1.400 1874.180 1279.600 ;
      RECT 1876.140 1.400 1876.420 1279.600 ;
      RECT 1878.380 1.400 1878.660 1279.600 ;
      RECT 1880.620 1.400 1880.900 1279.600 ;
      RECT 1882.860 1.400 1883.140 1279.600 ;
      RECT 1885.100 1.400 1885.380 1279.600 ;
      RECT 1887.340 1.400 1887.620 1279.600 ;
      RECT 1889.580 1.400 1889.860 1279.600 ;
      RECT 1891.820 1.400 1892.100 1279.600 ;
      RECT 1894.060 1.400 1894.340 1279.600 ;
      RECT 1896.300 1.400 1896.580 1279.600 ;
      RECT 1898.540 1.400 1898.820 1279.600 ;
      RECT 1900.780 1.400 1901.060 1279.600 ;
      RECT 1903.020 1.400 1903.300 1279.600 ;
      RECT 1905.260 1.400 1905.540 1279.600 ;
      RECT 1907.500 1.400 1907.780 1279.600 ;
      RECT 1909.740 1.400 1910.020 1279.600 ;
      RECT 1911.980 1.400 1912.260 1279.600 ;
      RECT 1914.220 1.400 1914.500 1279.600 ;
      RECT 1916.460 1.400 1916.740 1279.600 ;
      RECT 1918.700 1.400 1918.980 1279.600 ;
      RECT 1920.940 1.400 1921.220 1279.600 ;
      RECT 1923.180 1.400 1923.460 1279.600 ;
      RECT 1925.420 1.400 1925.700 1279.600 ;
      RECT 1927.660 1.400 1927.940 1279.600 ;
      RECT 1929.900 1.400 1930.180 1279.600 ;
      RECT 1932.140 1.400 1932.420 1279.600 ;
      RECT 1934.380 1.400 1934.660 1279.600 ;
      RECT 1936.620 1.400 1936.900 1279.600 ;
      RECT 1938.860 1.400 1939.140 1279.600 ;
      RECT 1941.100 1.400 1941.380 1279.600 ;
      RECT 1943.340 1.400 1943.620 1279.600 ;
      RECT 1945.580 1.400 1945.860 1279.600 ;
      RECT 1947.820 1.400 1948.100 1279.600 ;
      RECT 1950.060 1.400 1950.340 1279.600 ;
      RECT 1952.300 1.400 1952.580 1279.600 ;
      RECT 1954.540 1.400 1954.820 1279.600 ;
      RECT 1956.780 1.400 1957.060 1279.600 ;
      RECT 1959.020 1.400 1959.300 1279.600 ;
      RECT 1961.260 1.400 1961.540 1279.600 ;
      RECT 1963.500 1.400 1963.780 1279.600 ;
      RECT 1965.740 1.400 1966.020 1279.600 ;
      RECT 1967.980 1.400 1968.260 1279.600 ;
      RECT 1970.220 1.400 1970.500 1279.600 ;
      RECT 1972.460 1.400 1972.740 1279.600 ;
      RECT 1974.700 1.400 1974.980 1279.600 ;
      RECT 1976.940 1.400 1977.220 1279.600 ;
      RECT 1979.180 1.400 1979.460 1279.600 ;
      RECT 1981.420 1.400 1981.700 1279.600 ;
      RECT 1983.660 1.400 1983.940 1279.600 ;
      RECT 1985.900 1.400 1986.180 1279.600 ;
      RECT 1988.140 1.400 1988.420 1279.600 ;
      RECT 1990.380 1.400 1990.660 1279.600 ;
      RECT 1992.620 1.400 1992.900 1279.600 ;
      RECT 1994.860 1.400 1995.140 1279.600 ;
      RECT 1997.100 1.400 1997.380 1279.600 ;
      RECT 1999.340 1.400 1999.620 1279.600 ;
      RECT 2001.580 1.400 2001.860 1279.600 ;
      RECT 2003.820 1.400 2004.100 1279.600 ;
      RECT 2006.060 1.400 2006.340 1279.600 ;
      RECT 2008.300 1.400 2008.580 1279.600 ;
      RECT 2010.540 1.400 2010.820 1279.600 ;
      RECT 2012.780 1.400 2013.060 1279.600 ;
      RECT 2015.020 1.400 2015.300 1279.600 ;
      RECT 2017.260 1.400 2017.540 1279.600 ;
      RECT 2019.500 1.400 2019.780 1279.600 ;
      RECT 2021.740 1.400 2022.020 1279.600 ;
      RECT 2023.980 1.400 2024.260 1279.600 ;
      RECT 2026.220 1.400 2026.500 1279.600 ;
      RECT 2028.460 1.400 2028.740 1279.600 ;
      RECT 2030.700 1.400 2030.980 1279.600 ;
      RECT 2032.940 1.400 2033.220 1279.600 ;
      RECT 2035.180 1.400 2035.460 1279.600 ;
      RECT 2037.420 1.400 2037.700 1279.600 ;
      RECT 2039.660 1.400 2039.940 1279.600 ;
      RECT 2041.900 1.400 2042.180 1279.600 ;
      RECT 2044.140 1.400 2044.420 1279.600 ;
      RECT 2046.380 1.400 2046.660 1279.600 ;
      RECT 2048.620 1.400 2048.900 1279.600 ;
      RECT 2050.860 1.400 2051.140 1279.600 ;
      RECT 2053.100 1.400 2053.380 1279.600 ;
      RECT 2055.340 1.400 2055.620 1279.600 ;
      RECT 2057.580 1.400 2057.860 1279.600 ;
      RECT 2059.820 1.400 2060.100 1279.600 ;
      RECT 2062.060 1.400 2062.340 1279.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 1279.600 ;
      RECT 4.620 1.400 4.900 1279.600 ;
      RECT 6.860 1.400 7.140 1279.600 ;
      RECT 9.100 1.400 9.380 1279.600 ;
      RECT 11.340 1.400 11.620 1279.600 ;
      RECT 13.580 1.400 13.860 1279.600 ;
      RECT 15.820 1.400 16.100 1279.600 ;
      RECT 18.060 1.400 18.340 1279.600 ;
      RECT 20.300 1.400 20.580 1279.600 ;
      RECT 22.540 1.400 22.820 1279.600 ;
      RECT 24.780 1.400 25.060 1279.600 ;
      RECT 27.020 1.400 27.300 1279.600 ;
      RECT 29.260 1.400 29.540 1279.600 ;
      RECT 31.500 1.400 31.780 1279.600 ;
      RECT 33.740 1.400 34.020 1279.600 ;
      RECT 35.980 1.400 36.260 1279.600 ;
      RECT 38.220 1.400 38.500 1279.600 ;
      RECT 40.460 1.400 40.740 1279.600 ;
      RECT 42.700 1.400 42.980 1279.600 ;
      RECT 44.940 1.400 45.220 1279.600 ;
      RECT 47.180 1.400 47.460 1279.600 ;
      RECT 49.420 1.400 49.700 1279.600 ;
      RECT 51.660 1.400 51.940 1279.600 ;
      RECT 53.900 1.400 54.180 1279.600 ;
      RECT 56.140 1.400 56.420 1279.600 ;
      RECT 58.380 1.400 58.660 1279.600 ;
      RECT 60.620 1.400 60.900 1279.600 ;
      RECT 62.860 1.400 63.140 1279.600 ;
      RECT 65.100 1.400 65.380 1279.600 ;
      RECT 67.340 1.400 67.620 1279.600 ;
      RECT 69.580 1.400 69.860 1279.600 ;
      RECT 71.820 1.400 72.100 1279.600 ;
      RECT 74.060 1.400 74.340 1279.600 ;
      RECT 76.300 1.400 76.580 1279.600 ;
      RECT 78.540 1.400 78.820 1279.600 ;
      RECT 80.780 1.400 81.060 1279.600 ;
      RECT 83.020 1.400 83.300 1279.600 ;
      RECT 85.260 1.400 85.540 1279.600 ;
      RECT 87.500 1.400 87.780 1279.600 ;
      RECT 89.740 1.400 90.020 1279.600 ;
      RECT 91.980 1.400 92.260 1279.600 ;
      RECT 94.220 1.400 94.500 1279.600 ;
      RECT 96.460 1.400 96.740 1279.600 ;
      RECT 98.700 1.400 98.980 1279.600 ;
      RECT 100.940 1.400 101.220 1279.600 ;
      RECT 103.180 1.400 103.460 1279.600 ;
      RECT 105.420 1.400 105.700 1279.600 ;
      RECT 107.660 1.400 107.940 1279.600 ;
      RECT 109.900 1.400 110.180 1279.600 ;
      RECT 112.140 1.400 112.420 1279.600 ;
      RECT 114.380 1.400 114.660 1279.600 ;
      RECT 116.620 1.400 116.900 1279.600 ;
      RECT 118.860 1.400 119.140 1279.600 ;
      RECT 121.100 1.400 121.380 1279.600 ;
      RECT 123.340 1.400 123.620 1279.600 ;
      RECT 125.580 1.400 125.860 1279.600 ;
      RECT 127.820 1.400 128.100 1279.600 ;
      RECT 130.060 1.400 130.340 1279.600 ;
      RECT 132.300 1.400 132.580 1279.600 ;
      RECT 134.540 1.400 134.820 1279.600 ;
      RECT 136.780 1.400 137.060 1279.600 ;
      RECT 139.020 1.400 139.300 1279.600 ;
      RECT 141.260 1.400 141.540 1279.600 ;
      RECT 143.500 1.400 143.780 1279.600 ;
      RECT 145.740 1.400 146.020 1279.600 ;
      RECT 147.980 1.400 148.260 1279.600 ;
      RECT 150.220 1.400 150.500 1279.600 ;
      RECT 152.460 1.400 152.740 1279.600 ;
      RECT 154.700 1.400 154.980 1279.600 ;
      RECT 156.940 1.400 157.220 1279.600 ;
      RECT 159.180 1.400 159.460 1279.600 ;
      RECT 161.420 1.400 161.700 1279.600 ;
      RECT 163.660 1.400 163.940 1279.600 ;
      RECT 165.900 1.400 166.180 1279.600 ;
      RECT 168.140 1.400 168.420 1279.600 ;
      RECT 170.380 1.400 170.660 1279.600 ;
      RECT 172.620 1.400 172.900 1279.600 ;
      RECT 174.860 1.400 175.140 1279.600 ;
      RECT 177.100 1.400 177.380 1279.600 ;
      RECT 179.340 1.400 179.620 1279.600 ;
      RECT 181.580 1.400 181.860 1279.600 ;
      RECT 183.820 1.400 184.100 1279.600 ;
      RECT 186.060 1.400 186.340 1279.600 ;
      RECT 188.300 1.400 188.580 1279.600 ;
      RECT 190.540 1.400 190.820 1279.600 ;
      RECT 192.780 1.400 193.060 1279.600 ;
      RECT 195.020 1.400 195.300 1279.600 ;
      RECT 197.260 1.400 197.540 1279.600 ;
      RECT 199.500 1.400 199.780 1279.600 ;
      RECT 201.740 1.400 202.020 1279.600 ;
      RECT 203.980 1.400 204.260 1279.600 ;
      RECT 206.220 1.400 206.500 1279.600 ;
      RECT 208.460 1.400 208.740 1279.600 ;
      RECT 210.700 1.400 210.980 1279.600 ;
      RECT 212.940 1.400 213.220 1279.600 ;
      RECT 215.180 1.400 215.460 1279.600 ;
      RECT 217.420 1.400 217.700 1279.600 ;
      RECT 219.660 1.400 219.940 1279.600 ;
      RECT 221.900 1.400 222.180 1279.600 ;
      RECT 224.140 1.400 224.420 1279.600 ;
      RECT 226.380 1.400 226.660 1279.600 ;
      RECT 228.620 1.400 228.900 1279.600 ;
      RECT 230.860 1.400 231.140 1279.600 ;
      RECT 233.100 1.400 233.380 1279.600 ;
      RECT 235.340 1.400 235.620 1279.600 ;
      RECT 237.580 1.400 237.860 1279.600 ;
      RECT 239.820 1.400 240.100 1279.600 ;
      RECT 242.060 1.400 242.340 1279.600 ;
      RECT 244.300 1.400 244.580 1279.600 ;
      RECT 246.540 1.400 246.820 1279.600 ;
      RECT 248.780 1.400 249.060 1279.600 ;
      RECT 251.020 1.400 251.300 1279.600 ;
      RECT 253.260 1.400 253.540 1279.600 ;
      RECT 255.500 1.400 255.780 1279.600 ;
      RECT 257.740 1.400 258.020 1279.600 ;
      RECT 259.980 1.400 260.260 1279.600 ;
      RECT 262.220 1.400 262.500 1279.600 ;
      RECT 264.460 1.400 264.740 1279.600 ;
      RECT 266.700 1.400 266.980 1279.600 ;
      RECT 268.940 1.400 269.220 1279.600 ;
      RECT 271.180 1.400 271.460 1279.600 ;
      RECT 273.420 1.400 273.700 1279.600 ;
      RECT 275.660 1.400 275.940 1279.600 ;
      RECT 277.900 1.400 278.180 1279.600 ;
      RECT 280.140 1.400 280.420 1279.600 ;
      RECT 282.380 1.400 282.660 1279.600 ;
      RECT 284.620 1.400 284.900 1279.600 ;
      RECT 286.860 1.400 287.140 1279.600 ;
      RECT 289.100 1.400 289.380 1279.600 ;
      RECT 291.340 1.400 291.620 1279.600 ;
      RECT 293.580 1.400 293.860 1279.600 ;
      RECT 295.820 1.400 296.100 1279.600 ;
      RECT 298.060 1.400 298.340 1279.600 ;
      RECT 300.300 1.400 300.580 1279.600 ;
      RECT 302.540 1.400 302.820 1279.600 ;
      RECT 304.780 1.400 305.060 1279.600 ;
      RECT 307.020 1.400 307.300 1279.600 ;
      RECT 309.260 1.400 309.540 1279.600 ;
      RECT 311.500 1.400 311.780 1279.600 ;
      RECT 313.740 1.400 314.020 1279.600 ;
      RECT 315.980 1.400 316.260 1279.600 ;
      RECT 318.220 1.400 318.500 1279.600 ;
      RECT 320.460 1.400 320.740 1279.600 ;
      RECT 322.700 1.400 322.980 1279.600 ;
      RECT 324.940 1.400 325.220 1279.600 ;
      RECT 327.180 1.400 327.460 1279.600 ;
      RECT 329.420 1.400 329.700 1279.600 ;
      RECT 331.660 1.400 331.940 1279.600 ;
      RECT 333.900 1.400 334.180 1279.600 ;
      RECT 336.140 1.400 336.420 1279.600 ;
      RECT 338.380 1.400 338.660 1279.600 ;
      RECT 340.620 1.400 340.900 1279.600 ;
      RECT 342.860 1.400 343.140 1279.600 ;
      RECT 345.100 1.400 345.380 1279.600 ;
      RECT 347.340 1.400 347.620 1279.600 ;
      RECT 349.580 1.400 349.860 1279.600 ;
      RECT 351.820 1.400 352.100 1279.600 ;
      RECT 354.060 1.400 354.340 1279.600 ;
      RECT 356.300 1.400 356.580 1279.600 ;
      RECT 358.540 1.400 358.820 1279.600 ;
      RECT 360.780 1.400 361.060 1279.600 ;
      RECT 363.020 1.400 363.300 1279.600 ;
      RECT 365.260 1.400 365.540 1279.600 ;
      RECT 367.500 1.400 367.780 1279.600 ;
      RECT 369.740 1.400 370.020 1279.600 ;
      RECT 371.980 1.400 372.260 1279.600 ;
      RECT 374.220 1.400 374.500 1279.600 ;
      RECT 376.460 1.400 376.740 1279.600 ;
      RECT 378.700 1.400 378.980 1279.600 ;
      RECT 380.940 1.400 381.220 1279.600 ;
      RECT 383.180 1.400 383.460 1279.600 ;
      RECT 385.420 1.400 385.700 1279.600 ;
      RECT 387.660 1.400 387.940 1279.600 ;
      RECT 389.900 1.400 390.180 1279.600 ;
      RECT 392.140 1.400 392.420 1279.600 ;
      RECT 394.380 1.400 394.660 1279.600 ;
      RECT 396.620 1.400 396.900 1279.600 ;
      RECT 398.860 1.400 399.140 1279.600 ;
      RECT 401.100 1.400 401.380 1279.600 ;
      RECT 403.340 1.400 403.620 1279.600 ;
      RECT 405.580 1.400 405.860 1279.600 ;
      RECT 407.820 1.400 408.100 1279.600 ;
      RECT 410.060 1.400 410.340 1279.600 ;
      RECT 412.300 1.400 412.580 1279.600 ;
      RECT 414.540 1.400 414.820 1279.600 ;
      RECT 416.780 1.400 417.060 1279.600 ;
      RECT 419.020 1.400 419.300 1279.600 ;
      RECT 421.260 1.400 421.540 1279.600 ;
      RECT 423.500 1.400 423.780 1279.600 ;
      RECT 425.740 1.400 426.020 1279.600 ;
      RECT 427.980 1.400 428.260 1279.600 ;
      RECT 430.220 1.400 430.500 1279.600 ;
      RECT 432.460 1.400 432.740 1279.600 ;
      RECT 434.700 1.400 434.980 1279.600 ;
      RECT 436.940 1.400 437.220 1279.600 ;
      RECT 439.180 1.400 439.460 1279.600 ;
      RECT 441.420 1.400 441.700 1279.600 ;
      RECT 443.660 1.400 443.940 1279.600 ;
      RECT 445.900 1.400 446.180 1279.600 ;
      RECT 448.140 1.400 448.420 1279.600 ;
      RECT 450.380 1.400 450.660 1279.600 ;
      RECT 452.620 1.400 452.900 1279.600 ;
      RECT 454.860 1.400 455.140 1279.600 ;
      RECT 457.100 1.400 457.380 1279.600 ;
      RECT 459.340 1.400 459.620 1279.600 ;
      RECT 461.580 1.400 461.860 1279.600 ;
      RECT 463.820 1.400 464.100 1279.600 ;
      RECT 466.060 1.400 466.340 1279.600 ;
      RECT 468.300 1.400 468.580 1279.600 ;
      RECT 470.540 1.400 470.820 1279.600 ;
      RECT 472.780 1.400 473.060 1279.600 ;
      RECT 475.020 1.400 475.300 1279.600 ;
      RECT 477.260 1.400 477.540 1279.600 ;
      RECT 479.500 1.400 479.780 1279.600 ;
      RECT 481.740 1.400 482.020 1279.600 ;
      RECT 483.980 1.400 484.260 1279.600 ;
      RECT 486.220 1.400 486.500 1279.600 ;
      RECT 488.460 1.400 488.740 1279.600 ;
      RECT 490.700 1.400 490.980 1279.600 ;
      RECT 492.940 1.400 493.220 1279.600 ;
      RECT 495.180 1.400 495.460 1279.600 ;
      RECT 497.420 1.400 497.700 1279.600 ;
      RECT 499.660 1.400 499.940 1279.600 ;
      RECT 501.900 1.400 502.180 1279.600 ;
      RECT 504.140 1.400 504.420 1279.600 ;
      RECT 506.380 1.400 506.660 1279.600 ;
      RECT 508.620 1.400 508.900 1279.600 ;
      RECT 510.860 1.400 511.140 1279.600 ;
      RECT 513.100 1.400 513.380 1279.600 ;
      RECT 515.340 1.400 515.620 1279.600 ;
      RECT 517.580 1.400 517.860 1279.600 ;
      RECT 519.820 1.400 520.100 1279.600 ;
      RECT 522.060 1.400 522.340 1279.600 ;
      RECT 524.300 1.400 524.580 1279.600 ;
      RECT 526.540 1.400 526.820 1279.600 ;
      RECT 528.780 1.400 529.060 1279.600 ;
      RECT 531.020 1.400 531.300 1279.600 ;
      RECT 533.260 1.400 533.540 1279.600 ;
      RECT 535.500 1.400 535.780 1279.600 ;
      RECT 537.740 1.400 538.020 1279.600 ;
      RECT 539.980 1.400 540.260 1279.600 ;
      RECT 542.220 1.400 542.500 1279.600 ;
      RECT 544.460 1.400 544.740 1279.600 ;
      RECT 546.700 1.400 546.980 1279.600 ;
      RECT 548.940 1.400 549.220 1279.600 ;
      RECT 551.180 1.400 551.460 1279.600 ;
      RECT 553.420 1.400 553.700 1279.600 ;
      RECT 555.660 1.400 555.940 1279.600 ;
      RECT 557.900 1.400 558.180 1279.600 ;
      RECT 560.140 1.400 560.420 1279.600 ;
      RECT 562.380 1.400 562.660 1279.600 ;
      RECT 564.620 1.400 564.900 1279.600 ;
      RECT 566.860 1.400 567.140 1279.600 ;
      RECT 569.100 1.400 569.380 1279.600 ;
      RECT 571.340 1.400 571.620 1279.600 ;
      RECT 573.580 1.400 573.860 1279.600 ;
      RECT 575.820 1.400 576.100 1279.600 ;
      RECT 578.060 1.400 578.340 1279.600 ;
      RECT 580.300 1.400 580.580 1279.600 ;
      RECT 582.540 1.400 582.820 1279.600 ;
      RECT 584.780 1.400 585.060 1279.600 ;
      RECT 587.020 1.400 587.300 1279.600 ;
      RECT 589.260 1.400 589.540 1279.600 ;
      RECT 591.500 1.400 591.780 1279.600 ;
      RECT 593.740 1.400 594.020 1279.600 ;
      RECT 595.980 1.400 596.260 1279.600 ;
      RECT 598.220 1.400 598.500 1279.600 ;
      RECT 600.460 1.400 600.740 1279.600 ;
      RECT 602.700 1.400 602.980 1279.600 ;
      RECT 604.940 1.400 605.220 1279.600 ;
      RECT 607.180 1.400 607.460 1279.600 ;
      RECT 609.420 1.400 609.700 1279.600 ;
      RECT 611.660 1.400 611.940 1279.600 ;
      RECT 613.900 1.400 614.180 1279.600 ;
      RECT 616.140 1.400 616.420 1279.600 ;
      RECT 618.380 1.400 618.660 1279.600 ;
      RECT 620.620 1.400 620.900 1279.600 ;
      RECT 622.860 1.400 623.140 1279.600 ;
      RECT 625.100 1.400 625.380 1279.600 ;
      RECT 627.340 1.400 627.620 1279.600 ;
      RECT 629.580 1.400 629.860 1279.600 ;
      RECT 631.820 1.400 632.100 1279.600 ;
      RECT 634.060 1.400 634.340 1279.600 ;
      RECT 636.300 1.400 636.580 1279.600 ;
      RECT 638.540 1.400 638.820 1279.600 ;
      RECT 640.780 1.400 641.060 1279.600 ;
      RECT 643.020 1.400 643.300 1279.600 ;
      RECT 645.260 1.400 645.540 1279.600 ;
      RECT 647.500 1.400 647.780 1279.600 ;
      RECT 649.740 1.400 650.020 1279.600 ;
      RECT 651.980 1.400 652.260 1279.600 ;
      RECT 654.220 1.400 654.500 1279.600 ;
      RECT 656.460 1.400 656.740 1279.600 ;
      RECT 658.700 1.400 658.980 1279.600 ;
      RECT 660.940 1.400 661.220 1279.600 ;
      RECT 663.180 1.400 663.460 1279.600 ;
      RECT 665.420 1.400 665.700 1279.600 ;
      RECT 667.660 1.400 667.940 1279.600 ;
      RECT 669.900 1.400 670.180 1279.600 ;
      RECT 672.140 1.400 672.420 1279.600 ;
      RECT 674.380 1.400 674.660 1279.600 ;
      RECT 676.620 1.400 676.900 1279.600 ;
      RECT 678.860 1.400 679.140 1279.600 ;
      RECT 681.100 1.400 681.380 1279.600 ;
      RECT 683.340 1.400 683.620 1279.600 ;
      RECT 685.580 1.400 685.860 1279.600 ;
      RECT 687.820 1.400 688.100 1279.600 ;
      RECT 690.060 1.400 690.340 1279.600 ;
      RECT 692.300 1.400 692.580 1279.600 ;
      RECT 694.540 1.400 694.820 1279.600 ;
      RECT 696.780 1.400 697.060 1279.600 ;
      RECT 699.020 1.400 699.300 1279.600 ;
      RECT 701.260 1.400 701.540 1279.600 ;
      RECT 703.500 1.400 703.780 1279.600 ;
      RECT 705.740 1.400 706.020 1279.600 ;
      RECT 707.980 1.400 708.260 1279.600 ;
      RECT 710.220 1.400 710.500 1279.600 ;
      RECT 712.460 1.400 712.740 1279.600 ;
      RECT 714.700 1.400 714.980 1279.600 ;
      RECT 716.940 1.400 717.220 1279.600 ;
      RECT 719.180 1.400 719.460 1279.600 ;
      RECT 721.420 1.400 721.700 1279.600 ;
      RECT 723.660 1.400 723.940 1279.600 ;
      RECT 725.900 1.400 726.180 1279.600 ;
      RECT 728.140 1.400 728.420 1279.600 ;
      RECT 730.380 1.400 730.660 1279.600 ;
      RECT 732.620 1.400 732.900 1279.600 ;
      RECT 734.860 1.400 735.140 1279.600 ;
      RECT 737.100 1.400 737.380 1279.600 ;
      RECT 739.340 1.400 739.620 1279.600 ;
      RECT 741.580 1.400 741.860 1279.600 ;
      RECT 743.820 1.400 744.100 1279.600 ;
      RECT 746.060 1.400 746.340 1279.600 ;
      RECT 748.300 1.400 748.580 1279.600 ;
      RECT 750.540 1.400 750.820 1279.600 ;
      RECT 752.780 1.400 753.060 1279.600 ;
      RECT 755.020 1.400 755.300 1279.600 ;
      RECT 757.260 1.400 757.540 1279.600 ;
      RECT 759.500 1.400 759.780 1279.600 ;
      RECT 761.740 1.400 762.020 1279.600 ;
      RECT 763.980 1.400 764.260 1279.600 ;
      RECT 766.220 1.400 766.500 1279.600 ;
      RECT 768.460 1.400 768.740 1279.600 ;
      RECT 770.700 1.400 770.980 1279.600 ;
      RECT 772.940 1.400 773.220 1279.600 ;
      RECT 775.180 1.400 775.460 1279.600 ;
      RECT 777.420 1.400 777.700 1279.600 ;
      RECT 779.660 1.400 779.940 1279.600 ;
      RECT 781.900 1.400 782.180 1279.600 ;
      RECT 784.140 1.400 784.420 1279.600 ;
      RECT 786.380 1.400 786.660 1279.600 ;
      RECT 788.620 1.400 788.900 1279.600 ;
      RECT 790.860 1.400 791.140 1279.600 ;
      RECT 793.100 1.400 793.380 1279.600 ;
      RECT 795.340 1.400 795.620 1279.600 ;
      RECT 797.580 1.400 797.860 1279.600 ;
      RECT 799.820 1.400 800.100 1279.600 ;
      RECT 802.060 1.400 802.340 1279.600 ;
      RECT 804.300 1.400 804.580 1279.600 ;
      RECT 806.540 1.400 806.820 1279.600 ;
      RECT 808.780 1.400 809.060 1279.600 ;
      RECT 811.020 1.400 811.300 1279.600 ;
      RECT 813.260 1.400 813.540 1279.600 ;
      RECT 815.500 1.400 815.780 1279.600 ;
      RECT 817.740 1.400 818.020 1279.600 ;
      RECT 819.980 1.400 820.260 1279.600 ;
      RECT 822.220 1.400 822.500 1279.600 ;
      RECT 824.460 1.400 824.740 1279.600 ;
      RECT 826.700 1.400 826.980 1279.600 ;
      RECT 828.940 1.400 829.220 1279.600 ;
      RECT 831.180 1.400 831.460 1279.600 ;
      RECT 833.420 1.400 833.700 1279.600 ;
      RECT 835.660 1.400 835.940 1279.600 ;
      RECT 837.900 1.400 838.180 1279.600 ;
      RECT 840.140 1.400 840.420 1279.600 ;
      RECT 842.380 1.400 842.660 1279.600 ;
      RECT 844.620 1.400 844.900 1279.600 ;
      RECT 846.860 1.400 847.140 1279.600 ;
      RECT 849.100 1.400 849.380 1279.600 ;
      RECT 851.340 1.400 851.620 1279.600 ;
      RECT 853.580 1.400 853.860 1279.600 ;
      RECT 855.820 1.400 856.100 1279.600 ;
      RECT 858.060 1.400 858.340 1279.600 ;
      RECT 860.300 1.400 860.580 1279.600 ;
      RECT 862.540 1.400 862.820 1279.600 ;
      RECT 864.780 1.400 865.060 1279.600 ;
      RECT 867.020 1.400 867.300 1279.600 ;
      RECT 869.260 1.400 869.540 1279.600 ;
      RECT 871.500 1.400 871.780 1279.600 ;
      RECT 873.740 1.400 874.020 1279.600 ;
      RECT 875.980 1.400 876.260 1279.600 ;
      RECT 878.220 1.400 878.500 1279.600 ;
      RECT 880.460 1.400 880.740 1279.600 ;
      RECT 882.700 1.400 882.980 1279.600 ;
      RECT 884.940 1.400 885.220 1279.600 ;
      RECT 887.180 1.400 887.460 1279.600 ;
      RECT 889.420 1.400 889.700 1279.600 ;
      RECT 891.660 1.400 891.940 1279.600 ;
      RECT 893.900 1.400 894.180 1279.600 ;
      RECT 896.140 1.400 896.420 1279.600 ;
      RECT 898.380 1.400 898.660 1279.600 ;
      RECT 900.620 1.400 900.900 1279.600 ;
      RECT 902.860 1.400 903.140 1279.600 ;
      RECT 905.100 1.400 905.380 1279.600 ;
      RECT 907.340 1.400 907.620 1279.600 ;
      RECT 909.580 1.400 909.860 1279.600 ;
      RECT 911.820 1.400 912.100 1279.600 ;
      RECT 914.060 1.400 914.340 1279.600 ;
      RECT 916.300 1.400 916.580 1279.600 ;
      RECT 918.540 1.400 918.820 1279.600 ;
      RECT 920.780 1.400 921.060 1279.600 ;
      RECT 923.020 1.400 923.300 1279.600 ;
      RECT 925.260 1.400 925.540 1279.600 ;
      RECT 927.500 1.400 927.780 1279.600 ;
      RECT 929.740 1.400 930.020 1279.600 ;
      RECT 931.980 1.400 932.260 1279.600 ;
      RECT 934.220 1.400 934.500 1279.600 ;
      RECT 936.460 1.400 936.740 1279.600 ;
      RECT 938.700 1.400 938.980 1279.600 ;
      RECT 940.940 1.400 941.220 1279.600 ;
      RECT 943.180 1.400 943.460 1279.600 ;
      RECT 945.420 1.400 945.700 1279.600 ;
      RECT 947.660 1.400 947.940 1279.600 ;
      RECT 949.900 1.400 950.180 1279.600 ;
      RECT 952.140 1.400 952.420 1279.600 ;
      RECT 954.380 1.400 954.660 1279.600 ;
      RECT 956.620 1.400 956.900 1279.600 ;
      RECT 958.860 1.400 959.140 1279.600 ;
      RECT 961.100 1.400 961.380 1279.600 ;
      RECT 963.340 1.400 963.620 1279.600 ;
      RECT 965.580 1.400 965.860 1279.600 ;
      RECT 967.820 1.400 968.100 1279.600 ;
      RECT 970.060 1.400 970.340 1279.600 ;
      RECT 972.300 1.400 972.580 1279.600 ;
      RECT 974.540 1.400 974.820 1279.600 ;
      RECT 976.780 1.400 977.060 1279.600 ;
      RECT 979.020 1.400 979.300 1279.600 ;
      RECT 981.260 1.400 981.540 1279.600 ;
      RECT 983.500 1.400 983.780 1279.600 ;
      RECT 985.740 1.400 986.020 1279.600 ;
      RECT 987.980 1.400 988.260 1279.600 ;
      RECT 990.220 1.400 990.500 1279.600 ;
      RECT 992.460 1.400 992.740 1279.600 ;
      RECT 994.700 1.400 994.980 1279.600 ;
      RECT 996.940 1.400 997.220 1279.600 ;
      RECT 999.180 1.400 999.460 1279.600 ;
      RECT 1001.420 1.400 1001.700 1279.600 ;
      RECT 1003.660 1.400 1003.940 1279.600 ;
      RECT 1005.900 1.400 1006.180 1279.600 ;
      RECT 1008.140 1.400 1008.420 1279.600 ;
      RECT 1010.380 1.400 1010.660 1279.600 ;
      RECT 1012.620 1.400 1012.900 1279.600 ;
      RECT 1014.860 1.400 1015.140 1279.600 ;
      RECT 1017.100 1.400 1017.380 1279.600 ;
      RECT 1019.340 1.400 1019.620 1279.600 ;
      RECT 1021.580 1.400 1021.860 1279.600 ;
      RECT 1023.820 1.400 1024.100 1279.600 ;
      RECT 1026.060 1.400 1026.340 1279.600 ;
      RECT 1028.300 1.400 1028.580 1279.600 ;
      RECT 1030.540 1.400 1030.820 1279.600 ;
      RECT 1032.780 1.400 1033.060 1279.600 ;
      RECT 1035.020 1.400 1035.300 1279.600 ;
      RECT 1037.260 1.400 1037.540 1279.600 ;
      RECT 1039.500 1.400 1039.780 1279.600 ;
      RECT 1041.740 1.400 1042.020 1279.600 ;
      RECT 1043.980 1.400 1044.260 1279.600 ;
      RECT 1046.220 1.400 1046.500 1279.600 ;
      RECT 1048.460 1.400 1048.740 1279.600 ;
      RECT 1050.700 1.400 1050.980 1279.600 ;
      RECT 1052.940 1.400 1053.220 1279.600 ;
      RECT 1055.180 1.400 1055.460 1279.600 ;
      RECT 1057.420 1.400 1057.700 1279.600 ;
      RECT 1059.660 1.400 1059.940 1279.600 ;
      RECT 1061.900 1.400 1062.180 1279.600 ;
      RECT 1064.140 1.400 1064.420 1279.600 ;
      RECT 1066.380 1.400 1066.660 1279.600 ;
      RECT 1068.620 1.400 1068.900 1279.600 ;
      RECT 1070.860 1.400 1071.140 1279.600 ;
      RECT 1073.100 1.400 1073.380 1279.600 ;
      RECT 1075.340 1.400 1075.620 1279.600 ;
      RECT 1077.580 1.400 1077.860 1279.600 ;
      RECT 1079.820 1.400 1080.100 1279.600 ;
      RECT 1082.060 1.400 1082.340 1279.600 ;
      RECT 1084.300 1.400 1084.580 1279.600 ;
      RECT 1086.540 1.400 1086.820 1279.600 ;
      RECT 1088.780 1.400 1089.060 1279.600 ;
      RECT 1091.020 1.400 1091.300 1279.600 ;
      RECT 1093.260 1.400 1093.540 1279.600 ;
      RECT 1095.500 1.400 1095.780 1279.600 ;
      RECT 1097.740 1.400 1098.020 1279.600 ;
      RECT 1099.980 1.400 1100.260 1279.600 ;
      RECT 1102.220 1.400 1102.500 1279.600 ;
      RECT 1104.460 1.400 1104.740 1279.600 ;
      RECT 1106.700 1.400 1106.980 1279.600 ;
      RECT 1108.940 1.400 1109.220 1279.600 ;
      RECT 1111.180 1.400 1111.460 1279.600 ;
      RECT 1113.420 1.400 1113.700 1279.600 ;
      RECT 1115.660 1.400 1115.940 1279.600 ;
      RECT 1117.900 1.400 1118.180 1279.600 ;
      RECT 1120.140 1.400 1120.420 1279.600 ;
      RECT 1122.380 1.400 1122.660 1279.600 ;
      RECT 1124.620 1.400 1124.900 1279.600 ;
      RECT 1126.860 1.400 1127.140 1279.600 ;
      RECT 1129.100 1.400 1129.380 1279.600 ;
      RECT 1131.340 1.400 1131.620 1279.600 ;
      RECT 1133.580 1.400 1133.860 1279.600 ;
      RECT 1135.820 1.400 1136.100 1279.600 ;
      RECT 1138.060 1.400 1138.340 1279.600 ;
      RECT 1140.300 1.400 1140.580 1279.600 ;
      RECT 1142.540 1.400 1142.820 1279.600 ;
      RECT 1144.780 1.400 1145.060 1279.600 ;
      RECT 1147.020 1.400 1147.300 1279.600 ;
      RECT 1149.260 1.400 1149.540 1279.600 ;
      RECT 1151.500 1.400 1151.780 1279.600 ;
      RECT 1153.740 1.400 1154.020 1279.600 ;
      RECT 1155.980 1.400 1156.260 1279.600 ;
      RECT 1158.220 1.400 1158.500 1279.600 ;
      RECT 1160.460 1.400 1160.740 1279.600 ;
      RECT 1162.700 1.400 1162.980 1279.600 ;
      RECT 1164.940 1.400 1165.220 1279.600 ;
      RECT 1167.180 1.400 1167.460 1279.600 ;
      RECT 1169.420 1.400 1169.700 1279.600 ;
      RECT 1171.660 1.400 1171.940 1279.600 ;
      RECT 1173.900 1.400 1174.180 1279.600 ;
      RECT 1176.140 1.400 1176.420 1279.600 ;
      RECT 1178.380 1.400 1178.660 1279.600 ;
      RECT 1180.620 1.400 1180.900 1279.600 ;
      RECT 1182.860 1.400 1183.140 1279.600 ;
      RECT 1185.100 1.400 1185.380 1279.600 ;
      RECT 1187.340 1.400 1187.620 1279.600 ;
      RECT 1189.580 1.400 1189.860 1279.600 ;
      RECT 1191.820 1.400 1192.100 1279.600 ;
      RECT 1194.060 1.400 1194.340 1279.600 ;
      RECT 1196.300 1.400 1196.580 1279.600 ;
      RECT 1198.540 1.400 1198.820 1279.600 ;
      RECT 1200.780 1.400 1201.060 1279.600 ;
      RECT 1203.020 1.400 1203.300 1279.600 ;
      RECT 1205.260 1.400 1205.540 1279.600 ;
      RECT 1207.500 1.400 1207.780 1279.600 ;
      RECT 1209.740 1.400 1210.020 1279.600 ;
      RECT 1211.980 1.400 1212.260 1279.600 ;
      RECT 1214.220 1.400 1214.500 1279.600 ;
      RECT 1216.460 1.400 1216.740 1279.600 ;
      RECT 1218.700 1.400 1218.980 1279.600 ;
      RECT 1220.940 1.400 1221.220 1279.600 ;
      RECT 1223.180 1.400 1223.460 1279.600 ;
      RECT 1225.420 1.400 1225.700 1279.600 ;
      RECT 1227.660 1.400 1227.940 1279.600 ;
      RECT 1229.900 1.400 1230.180 1279.600 ;
      RECT 1232.140 1.400 1232.420 1279.600 ;
      RECT 1234.380 1.400 1234.660 1279.600 ;
      RECT 1236.620 1.400 1236.900 1279.600 ;
      RECT 1238.860 1.400 1239.140 1279.600 ;
      RECT 1241.100 1.400 1241.380 1279.600 ;
      RECT 1243.340 1.400 1243.620 1279.600 ;
      RECT 1245.580 1.400 1245.860 1279.600 ;
      RECT 1247.820 1.400 1248.100 1279.600 ;
      RECT 1250.060 1.400 1250.340 1279.600 ;
      RECT 1252.300 1.400 1252.580 1279.600 ;
      RECT 1254.540 1.400 1254.820 1279.600 ;
      RECT 1256.780 1.400 1257.060 1279.600 ;
      RECT 1259.020 1.400 1259.300 1279.600 ;
      RECT 1261.260 1.400 1261.540 1279.600 ;
      RECT 1263.500 1.400 1263.780 1279.600 ;
      RECT 1265.740 1.400 1266.020 1279.600 ;
      RECT 1267.980 1.400 1268.260 1279.600 ;
      RECT 1270.220 1.400 1270.500 1279.600 ;
      RECT 1272.460 1.400 1272.740 1279.600 ;
      RECT 1274.700 1.400 1274.980 1279.600 ;
      RECT 1276.940 1.400 1277.220 1279.600 ;
      RECT 1279.180 1.400 1279.460 1279.600 ;
      RECT 1281.420 1.400 1281.700 1279.600 ;
      RECT 1283.660 1.400 1283.940 1279.600 ;
      RECT 1285.900 1.400 1286.180 1279.600 ;
      RECT 1288.140 1.400 1288.420 1279.600 ;
      RECT 1290.380 1.400 1290.660 1279.600 ;
      RECT 1292.620 1.400 1292.900 1279.600 ;
      RECT 1294.860 1.400 1295.140 1279.600 ;
      RECT 1297.100 1.400 1297.380 1279.600 ;
      RECT 1299.340 1.400 1299.620 1279.600 ;
      RECT 1301.580 1.400 1301.860 1279.600 ;
      RECT 1303.820 1.400 1304.100 1279.600 ;
      RECT 1306.060 1.400 1306.340 1279.600 ;
      RECT 1308.300 1.400 1308.580 1279.600 ;
      RECT 1310.540 1.400 1310.820 1279.600 ;
      RECT 1312.780 1.400 1313.060 1279.600 ;
      RECT 1315.020 1.400 1315.300 1279.600 ;
      RECT 1317.260 1.400 1317.540 1279.600 ;
      RECT 1319.500 1.400 1319.780 1279.600 ;
      RECT 1321.740 1.400 1322.020 1279.600 ;
      RECT 1323.980 1.400 1324.260 1279.600 ;
      RECT 1326.220 1.400 1326.500 1279.600 ;
      RECT 1328.460 1.400 1328.740 1279.600 ;
      RECT 1330.700 1.400 1330.980 1279.600 ;
      RECT 1332.940 1.400 1333.220 1279.600 ;
      RECT 1335.180 1.400 1335.460 1279.600 ;
      RECT 1337.420 1.400 1337.700 1279.600 ;
      RECT 1339.660 1.400 1339.940 1279.600 ;
      RECT 1341.900 1.400 1342.180 1279.600 ;
      RECT 1344.140 1.400 1344.420 1279.600 ;
      RECT 1346.380 1.400 1346.660 1279.600 ;
      RECT 1348.620 1.400 1348.900 1279.600 ;
      RECT 1350.860 1.400 1351.140 1279.600 ;
      RECT 1353.100 1.400 1353.380 1279.600 ;
      RECT 1355.340 1.400 1355.620 1279.600 ;
      RECT 1357.580 1.400 1357.860 1279.600 ;
      RECT 1359.820 1.400 1360.100 1279.600 ;
      RECT 1362.060 1.400 1362.340 1279.600 ;
      RECT 1364.300 1.400 1364.580 1279.600 ;
      RECT 1366.540 1.400 1366.820 1279.600 ;
      RECT 1368.780 1.400 1369.060 1279.600 ;
      RECT 1371.020 1.400 1371.300 1279.600 ;
      RECT 1373.260 1.400 1373.540 1279.600 ;
      RECT 1375.500 1.400 1375.780 1279.600 ;
      RECT 1377.740 1.400 1378.020 1279.600 ;
      RECT 1379.980 1.400 1380.260 1279.600 ;
      RECT 1382.220 1.400 1382.500 1279.600 ;
      RECT 1384.460 1.400 1384.740 1279.600 ;
      RECT 1386.700 1.400 1386.980 1279.600 ;
      RECT 1388.940 1.400 1389.220 1279.600 ;
      RECT 1391.180 1.400 1391.460 1279.600 ;
      RECT 1393.420 1.400 1393.700 1279.600 ;
      RECT 1395.660 1.400 1395.940 1279.600 ;
      RECT 1397.900 1.400 1398.180 1279.600 ;
      RECT 1400.140 1.400 1400.420 1279.600 ;
      RECT 1402.380 1.400 1402.660 1279.600 ;
      RECT 1404.620 1.400 1404.900 1279.600 ;
      RECT 1406.860 1.400 1407.140 1279.600 ;
      RECT 1409.100 1.400 1409.380 1279.600 ;
      RECT 1411.340 1.400 1411.620 1279.600 ;
      RECT 1413.580 1.400 1413.860 1279.600 ;
      RECT 1415.820 1.400 1416.100 1279.600 ;
      RECT 1418.060 1.400 1418.340 1279.600 ;
      RECT 1420.300 1.400 1420.580 1279.600 ;
      RECT 1422.540 1.400 1422.820 1279.600 ;
      RECT 1424.780 1.400 1425.060 1279.600 ;
      RECT 1427.020 1.400 1427.300 1279.600 ;
      RECT 1429.260 1.400 1429.540 1279.600 ;
      RECT 1431.500 1.400 1431.780 1279.600 ;
      RECT 1433.740 1.400 1434.020 1279.600 ;
      RECT 1435.980 1.400 1436.260 1279.600 ;
      RECT 1438.220 1.400 1438.500 1279.600 ;
      RECT 1440.460 1.400 1440.740 1279.600 ;
      RECT 1442.700 1.400 1442.980 1279.600 ;
      RECT 1444.940 1.400 1445.220 1279.600 ;
      RECT 1447.180 1.400 1447.460 1279.600 ;
      RECT 1449.420 1.400 1449.700 1279.600 ;
      RECT 1451.660 1.400 1451.940 1279.600 ;
      RECT 1453.900 1.400 1454.180 1279.600 ;
      RECT 1456.140 1.400 1456.420 1279.600 ;
      RECT 1458.380 1.400 1458.660 1279.600 ;
      RECT 1460.620 1.400 1460.900 1279.600 ;
      RECT 1462.860 1.400 1463.140 1279.600 ;
      RECT 1465.100 1.400 1465.380 1279.600 ;
      RECT 1467.340 1.400 1467.620 1279.600 ;
      RECT 1469.580 1.400 1469.860 1279.600 ;
      RECT 1471.820 1.400 1472.100 1279.600 ;
      RECT 1474.060 1.400 1474.340 1279.600 ;
      RECT 1476.300 1.400 1476.580 1279.600 ;
      RECT 1478.540 1.400 1478.820 1279.600 ;
      RECT 1480.780 1.400 1481.060 1279.600 ;
      RECT 1483.020 1.400 1483.300 1279.600 ;
      RECT 1485.260 1.400 1485.540 1279.600 ;
      RECT 1487.500 1.400 1487.780 1279.600 ;
      RECT 1489.740 1.400 1490.020 1279.600 ;
      RECT 1491.980 1.400 1492.260 1279.600 ;
      RECT 1494.220 1.400 1494.500 1279.600 ;
      RECT 1496.460 1.400 1496.740 1279.600 ;
      RECT 1498.700 1.400 1498.980 1279.600 ;
      RECT 1500.940 1.400 1501.220 1279.600 ;
      RECT 1503.180 1.400 1503.460 1279.600 ;
      RECT 1505.420 1.400 1505.700 1279.600 ;
      RECT 1507.660 1.400 1507.940 1279.600 ;
      RECT 1509.900 1.400 1510.180 1279.600 ;
      RECT 1512.140 1.400 1512.420 1279.600 ;
      RECT 1514.380 1.400 1514.660 1279.600 ;
      RECT 1516.620 1.400 1516.900 1279.600 ;
      RECT 1518.860 1.400 1519.140 1279.600 ;
      RECT 1521.100 1.400 1521.380 1279.600 ;
      RECT 1523.340 1.400 1523.620 1279.600 ;
      RECT 1525.580 1.400 1525.860 1279.600 ;
      RECT 1527.820 1.400 1528.100 1279.600 ;
      RECT 1530.060 1.400 1530.340 1279.600 ;
      RECT 1532.300 1.400 1532.580 1279.600 ;
      RECT 1534.540 1.400 1534.820 1279.600 ;
      RECT 1536.780 1.400 1537.060 1279.600 ;
      RECT 1539.020 1.400 1539.300 1279.600 ;
      RECT 1541.260 1.400 1541.540 1279.600 ;
      RECT 1543.500 1.400 1543.780 1279.600 ;
      RECT 1545.740 1.400 1546.020 1279.600 ;
      RECT 1547.980 1.400 1548.260 1279.600 ;
      RECT 1550.220 1.400 1550.500 1279.600 ;
      RECT 1552.460 1.400 1552.740 1279.600 ;
      RECT 1554.700 1.400 1554.980 1279.600 ;
      RECT 1556.940 1.400 1557.220 1279.600 ;
      RECT 1559.180 1.400 1559.460 1279.600 ;
      RECT 1561.420 1.400 1561.700 1279.600 ;
      RECT 1563.660 1.400 1563.940 1279.600 ;
      RECT 1565.900 1.400 1566.180 1279.600 ;
      RECT 1568.140 1.400 1568.420 1279.600 ;
      RECT 1570.380 1.400 1570.660 1279.600 ;
      RECT 1572.620 1.400 1572.900 1279.600 ;
      RECT 1574.860 1.400 1575.140 1279.600 ;
      RECT 1577.100 1.400 1577.380 1279.600 ;
      RECT 1579.340 1.400 1579.620 1279.600 ;
      RECT 1581.580 1.400 1581.860 1279.600 ;
      RECT 1583.820 1.400 1584.100 1279.600 ;
      RECT 1586.060 1.400 1586.340 1279.600 ;
      RECT 1588.300 1.400 1588.580 1279.600 ;
      RECT 1590.540 1.400 1590.820 1279.600 ;
      RECT 1592.780 1.400 1593.060 1279.600 ;
      RECT 1595.020 1.400 1595.300 1279.600 ;
      RECT 1597.260 1.400 1597.540 1279.600 ;
      RECT 1599.500 1.400 1599.780 1279.600 ;
      RECT 1601.740 1.400 1602.020 1279.600 ;
      RECT 1603.980 1.400 1604.260 1279.600 ;
      RECT 1606.220 1.400 1606.500 1279.600 ;
      RECT 1608.460 1.400 1608.740 1279.600 ;
      RECT 1610.700 1.400 1610.980 1279.600 ;
      RECT 1612.940 1.400 1613.220 1279.600 ;
      RECT 1615.180 1.400 1615.460 1279.600 ;
      RECT 1617.420 1.400 1617.700 1279.600 ;
      RECT 1619.660 1.400 1619.940 1279.600 ;
      RECT 1621.900 1.400 1622.180 1279.600 ;
      RECT 1624.140 1.400 1624.420 1279.600 ;
      RECT 1626.380 1.400 1626.660 1279.600 ;
      RECT 1628.620 1.400 1628.900 1279.600 ;
      RECT 1630.860 1.400 1631.140 1279.600 ;
      RECT 1633.100 1.400 1633.380 1279.600 ;
      RECT 1635.340 1.400 1635.620 1279.600 ;
      RECT 1637.580 1.400 1637.860 1279.600 ;
      RECT 1639.820 1.400 1640.100 1279.600 ;
      RECT 1642.060 1.400 1642.340 1279.600 ;
      RECT 1644.300 1.400 1644.580 1279.600 ;
      RECT 1646.540 1.400 1646.820 1279.600 ;
      RECT 1648.780 1.400 1649.060 1279.600 ;
      RECT 1651.020 1.400 1651.300 1279.600 ;
      RECT 1653.260 1.400 1653.540 1279.600 ;
      RECT 1655.500 1.400 1655.780 1279.600 ;
      RECT 1657.740 1.400 1658.020 1279.600 ;
      RECT 1659.980 1.400 1660.260 1279.600 ;
      RECT 1662.220 1.400 1662.500 1279.600 ;
      RECT 1664.460 1.400 1664.740 1279.600 ;
      RECT 1666.700 1.400 1666.980 1279.600 ;
      RECT 1668.940 1.400 1669.220 1279.600 ;
      RECT 1671.180 1.400 1671.460 1279.600 ;
      RECT 1673.420 1.400 1673.700 1279.600 ;
      RECT 1675.660 1.400 1675.940 1279.600 ;
      RECT 1677.900 1.400 1678.180 1279.600 ;
      RECT 1680.140 1.400 1680.420 1279.600 ;
      RECT 1682.380 1.400 1682.660 1279.600 ;
      RECT 1684.620 1.400 1684.900 1279.600 ;
      RECT 1686.860 1.400 1687.140 1279.600 ;
      RECT 1689.100 1.400 1689.380 1279.600 ;
      RECT 1691.340 1.400 1691.620 1279.600 ;
      RECT 1693.580 1.400 1693.860 1279.600 ;
      RECT 1695.820 1.400 1696.100 1279.600 ;
      RECT 1698.060 1.400 1698.340 1279.600 ;
      RECT 1700.300 1.400 1700.580 1279.600 ;
      RECT 1702.540 1.400 1702.820 1279.600 ;
      RECT 1704.780 1.400 1705.060 1279.600 ;
      RECT 1707.020 1.400 1707.300 1279.600 ;
      RECT 1709.260 1.400 1709.540 1279.600 ;
      RECT 1711.500 1.400 1711.780 1279.600 ;
      RECT 1713.740 1.400 1714.020 1279.600 ;
      RECT 1715.980 1.400 1716.260 1279.600 ;
      RECT 1718.220 1.400 1718.500 1279.600 ;
      RECT 1720.460 1.400 1720.740 1279.600 ;
      RECT 1722.700 1.400 1722.980 1279.600 ;
      RECT 1724.940 1.400 1725.220 1279.600 ;
      RECT 1727.180 1.400 1727.460 1279.600 ;
      RECT 1729.420 1.400 1729.700 1279.600 ;
      RECT 1731.660 1.400 1731.940 1279.600 ;
      RECT 1733.900 1.400 1734.180 1279.600 ;
      RECT 1736.140 1.400 1736.420 1279.600 ;
      RECT 1738.380 1.400 1738.660 1279.600 ;
      RECT 1740.620 1.400 1740.900 1279.600 ;
      RECT 1742.860 1.400 1743.140 1279.600 ;
      RECT 1745.100 1.400 1745.380 1279.600 ;
      RECT 1747.340 1.400 1747.620 1279.600 ;
      RECT 1749.580 1.400 1749.860 1279.600 ;
      RECT 1751.820 1.400 1752.100 1279.600 ;
      RECT 1754.060 1.400 1754.340 1279.600 ;
      RECT 1756.300 1.400 1756.580 1279.600 ;
      RECT 1758.540 1.400 1758.820 1279.600 ;
      RECT 1760.780 1.400 1761.060 1279.600 ;
      RECT 1763.020 1.400 1763.300 1279.600 ;
      RECT 1765.260 1.400 1765.540 1279.600 ;
      RECT 1767.500 1.400 1767.780 1279.600 ;
      RECT 1769.740 1.400 1770.020 1279.600 ;
      RECT 1771.980 1.400 1772.260 1279.600 ;
      RECT 1774.220 1.400 1774.500 1279.600 ;
      RECT 1776.460 1.400 1776.740 1279.600 ;
      RECT 1778.700 1.400 1778.980 1279.600 ;
      RECT 1780.940 1.400 1781.220 1279.600 ;
      RECT 1783.180 1.400 1783.460 1279.600 ;
      RECT 1785.420 1.400 1785.700 1279.600 ;
      RECT 1787.660 1.400 1787.940 1279.600 ;
      RECT 1789.900 1.400 1790.180 1279.600 ;
      RECT 1792.140 1.400 1792.420 1279.600 ;
      RECT 1794.380 1.400 1794.660 1279.600 ;
      RECT 1796.620 1.400 1796.900 1279.600 ;
      RECT 1798.860 1.400 1799.140 1279.600 ;
      RECT 1801.100 1.400 1801.380 1279.600 ;
      RECT 1803.340 1.400 1803.620 1279.600 ;
      RECT 1805.580 1.400 1805.860 1279.600 ;
      RECT 1807.820 1.400 1808.100 1279.600 ;
      RECT 1810.060 1.400 1810.340 1279.600 ;
      RECT 1812.300 1.400 1812.580 1279.600 ;
      RECT 1814.540 1.400 1814.820 1279.600 ;
      RECT 1816.780 1.400 1817.060 1279.600 ;
      RECT 1819.020 1.400 1819.300 1279.600 ;
      RECT 1821.260 1.400 1821.540 1279.600 ;
      RECT 1823.500 1.400 1823.780 1279.600 ;
      RECT 1825.740 1.400 1826.020 1279.600 ;
      RECT 1827.980 1.400 1828.260 1279.600 ;
      RECT 1830.220 1.400 1830.500 1279.600 ;
      RECT 1832.460 1.400 1832.740 1279.600 ;
      RECT 1834.700 1.400 1834.980 1279.600 ;
      RECT 1836.940 1.400 1837.220 1279.600 ;
      RECT 1839.180 1.400 1839.460 1279.600 ;
      RECT 1841.420 1.400 1841.700 1279.600 ;
      RECT 1843.660 1.400 1843.940 1279.600 ;
      RECT 1845.900 1.400 1846.180 1279.600 ;
      RECT 1848.140 1.400 1848.420 1279.600 ;
      RECT 1850.380 1.400 1850.660 1279.600 ;
      RECT 1852.620 1.400 1852.900 1279.600 ;
      RECT 1854.860 1.400 1855.140 1279.600 ;
      RECT 1857.100 1.400 1857.380 1279.600 ;
      RECT 1859.340 1.400 1859.620 1279.600 ;
      RECT 1861.580 1.400 1861.860 1279.600 ;
      RECT 1863.820 1.400 1864.100 1279.600 ;
      RECT 1866.060 1.400 1866.340 1279.600 ;
      RECT 1868.300 1.400 1868.580 1279.600 ;
      RECT 1870.540 1.400 1870.820 1279.600 ;
      RECT 1872.780 1.400 1873.060 1279.600 ;
      RECT 1875.020 1.400 1875.300 1279.600 ;
      RECT 1877.260 1.400 1877.540 1279.600 ;
      RECT 1879.500 1.400 1879.780 1279.600 ;
      RECT 1881.740 1.400 1882.020 1279.600 ;
      RECT 1883.980 1.400 1884.260 1279.600 ;
      RECT 1886.220 1.400 1886.500 1279.600 ;
      RECT 1888.460 1.400 1888.740 1279.600 ;
      RECT 1890.700 1.400 1890.980 1279.600 ;
      RECT 1892.940 1.400 1893.220 1279.600 ;
      RECT 1895.180 1.400 1895.460 1279.600 ;
      RECT 1897.420 1.400 1897.700 1279.600 ;
      RECT 1899.660 1.400 1899.940 1279.600 ;
      RECT 1901.900 1.400 1902.180 1279.600 ;
      RECT 1904.140 1.400 1904.420 1279.600 ;
      RECT 1906.380 1.400 1906.660 1279.600 ;
      RECT 1908.620 1.400 1908.900 1279.600 ;
      RECT 1910.860 1.400 1911.140 1279.600 ;
      RECT 1913.100 1.400 1913.380 1279.600 ;
      RECT 1915.340 1.400 1915.620 1279.600 ;
      RECT 1917.580 1.400 1917.860 1279.600 ;
      RECT 1919.820 1.400 1920.100 1279.600 ;
      RECT 1922.060 1.400 1922.340 1279.600 ;
      RECT 1924.300 1.400 1924.580 1279.600 ;
      RECT 1926.540 1.400 1926.820 1279.600 ;
      RECT 1928.780 1.400 1929.060 1279.600 ;
      RECT 1931.020 1.400 1931.300 1279.600 ;
      RECT 1933.260 1.400 1933.540 1279.600 ;
      RECT 1935.500 1.400 1935.780 1279.600 ;
      RECT 1937.740 1.400 1938.020 1279.600 ;
      RECT 1939.980 1.400 1940.260 1279.600 ;
      RECT 1942.220 1.400 1942.500 1279.600 ;
      RECT 1944.460 1.400 1944.740 1279.600 ;
      RECT 1946.700 1.400 1946.980 1279.600 ;
      RECT 1948.940 1.400 1949.220 1279.600 ;
      RECT 1951.180 1.400 1951.460 1279.600 ;
      RECT 1953.420 1.400 1953.700 1279.600 ;
      RECT 1955.660 1.400 1955.940 1279.600 ;
      RECT 1957.900 1.400 1958.180 1279.600 ;
      RECT 1960.140 1.400 1960.420 1279.600 ;
      RECT 1962.380 1.400 1962.660 1279.600 ;
      RECT 1964.620 1.400 1964.900 1279.600 ;
      RECT 1966.860 1.400 1967.140 1279.600 ;
      RECT 1969.100 1.400 1969.380 1279.600 ;
      RECT 1971.340 1.400 1971.620 1279.600 ;
      RECT 1973.580 1.400 1973.860 1279.600 ;
      RECT 1975.820 1.400 1976.100 1279.600 ;
      RECT 1978.060 1.400 1978.340 1279.600 ;
      RECT 1980.300 1.400 1980.580 1279.600 ;
      RECT 1982.540 1.400 1982.820 1279.600 ;
      RECT 1984.780 1.400 1985.060 1279.600 ;
      RECT 1987.020 1.400 1987.300 1279.600 ;
      RECT 1989.260 1.400 1989.540 1279.600 ;
      RECT 1991.500 1.400 1991.780 1279.600 ;
      RECT 1993.740 1.400 1994.020 1279.600 ;
      RECT 1995.980 1.400 1996.260 1279.600 ;
      RECT 1998.220 1.400 1998.500 1279.600 ;
      RECT 2000.460 1.400 2000.740 1279.600 ;
      RECT 2002.700 1.400 2002.980 1279.600 ;
      RECT 2004.940 1.400 2005.220 1279.600 ;
      RECT 2007.180 1.400 2007.460 1279.600 ;
      RECT 2009.420 1.400 2009.700 1279.600 ;
      RECT 2011.660 1.400 2011.940 1279.600 ;
      RECT 2013.900 1.400 2014.180 1279.600 ;
      RECT 2016.140 1.400 2016.420 1279.600 ;
      RECT 2018.380 1.400 2018.660 1279.600 ;
      RECT 2020.620 1.400 2020.900 1279.600 ;
      RECT 2022.860 1.400 2023.140 1279.600 ;
      RECT 2025.100 1.400 2025.380 1279.600 ;
      RECT 2027.340 1.400 2027.620 1279.600 ;
      RECT 2029.580 1.400 2029.860 1279.600 ;
      RECT 2031.820 1.400 2032.100 1279.600 ;
      RECT 2034.060 1.400 2034.340 1279.600 ;
      RECT 2036.300 1.400 2036.580 1279.600 ;
      RECT 2038.540 1.400 2038.820 1279.600 ;
      RECT 2040.780 1.400 2041.060 1279.600 ;
      RECT 2043.020 1.400 2043.300 1279.600 ;
      RECT 2045.260 1.400 2045.540 1279.600 ;
      RECT 2047.500 1.400 2047.780 1279.600 ;
      RECT 2049.740 1.400 2050.020 1279.600 ;
      RECT 2051.980 1.400 2052.260 1279.600 ;
      RECT 2054.220 1.400 2054.500 1279.600 ;
      RECT 2056.460 1.400 2056.740 1279.600 ;
      RECT 2058.700 1.400 2058.980 1279.600 ;
      RECT 2060.940 1.400 2061.220 1279.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 2064.540 1281.000 ;
    LAYER metal2 ;
    RECT 0 0 2064.540 1281.000 ;
    LAYER metal3 ;
    RECT 0.070 0 2064.540 1281.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.065 ;
    RECT 0 2.135 0.070 2.765 ;
    RECT 0 2.835 0.070 3.465 ;
    RECT 0 3.535 0.070 4.165 ;
    RECT 0 4.235 0.070 4.865 ;
    RECT 0 4.935 0.070 5.565 ;
    RECT 0 5.635 0.070 6.265 ;
    RECT 0 6.335 0.070 6.965 ;
    RECT 0 7.035 0.070 7.665 ;
    RECT 0 7.735 0.070 8.365 ;
    RECT 0 8.435 0.070 9.065 ;
    RECT 0 9.135 0.070 9.765 ;
    RECT 0 9.835 0.070 10.465 ;
    RECT 0 10.535 0.070 11.165 ;
    RECT 0 11.235 0.070 11.865 ;
    RECT 0 11.935 0.070 12.565 ;
    RECT 0 12.635 0.070 13.265 ;
    RECT 0 13.335 0.070 13.965 ;
    RECT 0 14.035 0.070 14.665 ;
    RECT 0 14.735 0.070 15.365 ;
    RECT 0 15.435 0.070 16.065 ;
    RECT 0 16.135 0.070 16.765 ;
    RECT 0 16.835 0.070 17.465 ;
    RECT 0 17.535 0.070 18.165 ;
    RECT 0 18.235 0.070 18.865 ;
    RECT 0 18.935 0.070 19.565 ;
    RECT 0 19.635 0.070 20.265 ;
    RECT 0 20.335 0.070 20.965 ;
    RECT 0 21.035 0.070 21.665 ;
    RECT 0 21.735 0.070 22.365 ;
    RECT 0 22.435 0.070 23.065 ;
    RECT 0 23.135 0.070 23.765 ;
    RECT 0 23.835 0.070 24.465 ;
    RECT 0 24.535 0.070 25.165 ;
    RECT 0 25.235 0.070 25.865 ;
    RECT 0 25.935 0.070 26.565 ;
    RECT 0 26.635 0.070 27.265 ;
    RECT 0 27.335 0.070 27.965 ;
    RECT 0 28.035 0.070 28.665 ;
    RECT 0 28.735 0.070 29.365 ;
    RECT 0 29.435 0.070 30.065 ;
    RECT 0 30.135 0.070 30.765 ;
    RECT 0 30.835 0.070 31.465 ;
    RECT 0 31.535 0.070 32.165 ;
    RECT 0 32.235 0.070 32.865 ;
    RECT 0 32.935 0.070 33.565 ;
    RECT 0 33.635 0.070 34.265 ;
    RECT 0 34.335 0.070 34.965 ;
    RECT 0 35.035 0.070 35.665 ;
    RECT 0 35.735 0.070 36.365 ;
    RECT 0 36.435 0.070 37.065 ;
    RECT 0 37.135 0.070 37.765 ;
    RECT 0 37.835 0.070 38.465 ;
    RECT 0 38.535 0.070 39.165 ;
    RECT 0 39.235 0.070 39.865 ;
    RECT 0 39.935 0.070 40.565 ;
    RECT 0 40.635 0.070 41.265 ;
    RECT 0 41.335 0.070 41.965 ;
    RECT 0 42.035 0.070 42.665 ;
    RECT 0 42.735 0.070 43.365 ;
    RECT 0 43.435 0.070 44.065 ;
    RECT 0 44.135 0.070 44.765 ;
    RECT 0 44.835 0.070 45.465 ;
    RECT 0 45.535 0.070 46.165 ;
    RECT 0 46.235 0.070 46.865 ;
    RECT 0 46.935 0.070 47.565 ;
    RECT 0 47.635 0.070 48.265 ;
    RECT 0 48.335 0.070 48.965 ;
    RECT 0 49.035 0.070 49.665 ;
    RECT 0 49.735 0.070 50.365 ;
    RECT 0 50.435 0.070 51.065 ;
    RECT 0 51.135 0.070 51.765 ;
    RECT 0 51.835 0.070 52.465 ;
    RECT 0 52.535 0.070 53.165 ;
    RECT 0 53.235 0.070 53.865 ;
    RECT 0 53.935 0.070 54.565 ;
    RECT 0 54.635 0.070 55.265 ;
    RECT 0 55.335 0.070 55.965 ;
    RECT 0 56.035 0.070 56.665 ;
    RECT 0 56.735 0.070 57.365 ;
    RECT 0 57.435 0.070 58.065 ;
    RECT 0 58.135 0.070 58.765 ;
    RECT 0 58.835 0.070 59.465 ;
    RECT 0 59.535 0.070 60.165 ;
    RECT 0 60.235 0.070 60.865 ;
    RECT 0 60.935 0.070 61.565 ;
    RECT 0 61.635 0.070 62.265 ;
    RECT 0 62.335 0.070 62.965 ;
    RECT 0 63.035 0.070 63.665 ;
    RECT 0 63.735 0.070 64.365 ;
    RECT 0 64.435 0.070 65.065 ;
    RECT 0 65.135 0.070 65.765 ;
    RECT 0 65.835 0.070 66.465 ;
    RECT 0 66.535 0.070 67.165 ;
    RECT 0 67.235 0.070 67.865 ;
    RECT 0 67.935 0.070 68.565 ;
    RECT 0 68.635 0.070 69.265 ;
    RECT 0 69.335 0.070 69.965 ;
    RECT 0 70.035 0.070 70.665 ;
    RECT 0 70.735 0.070 71.365 ;
    RECT 0 71.435 0.070 72.065 ;
    RECT 0 72.135 0.070 72.765 ;
    RECT 0 72.835 0.070 73.465 ;
    RECT 0 73.535 0.070 74.165 ;
    RECT 0 74.235 0.070 74.865 ;
    RECT 0 74.935 0.070 75.565 ;
    RECT 0 75.635 0.070 76.265 ;
    RECT 0 76.335 0.070 76.965 ;
    RECT 0 77.035 0.070 77.665 ;
    RECT 0 77.735 0.070 78.365 ;
    RECT 0 78.435 0.070 79.065 ;
    RECT 0 79.135 0.070 79.765 ;
    RECT 0 79.835 0.070 80.465 ;
    RECT 0 80.535 0.070 81.165 ;
    RECT 0 81.235 0.070 81.865 ;
    RECT 0 81.935 0.070 82.565 ;
    RECT 0 82.635 0.070 83.265 ;
    RECT 0 83.335 0.070 83.965 ;
    RECT 0 84.035 0.070 84.665 ;
    RECT 0 84.735 0.070 85.365 ;
    RECT 0 85.435 0.070 86.065 ;
    RECT 0 86.135 0.070 86.765 ;
    RECT 0 86.835 0.070 87.465 ;
    RECT 0 87.535 0.070 88.165 ;
    RECT 0 88.235 0.070 88.865 ;
    RECT 0 88.935 0.070 89.565 ;
    RECT 0 89.635 0.070 90.265 ;
    RECT 0 90.335 0.070 90.965 ;
    RECT 0 91.035 0.070 91.665 ;
    RECT 0 91.735 0.070 92.365 ;
    RECT 0 92.435 0.070 93.065 ;
    RECT 0 93.135 0.070 93.765 ;
    RECT 0 93.835 0.070 94.465 ;
    RECT 0 94.535 0.070 95.165 ;
    RECT 0 95.235 0.070 95.865 ;
    RECT 0 95.935 0.070 96.565 ;
    RECT 0 96.635 0.070 97.265 ;
    RECT 0 97.335 0.070 97.965 ;
    RECT 0 98.035 0.070 98.665 ;
    RECT 0 98.735 0.070 99.365 ;
    RECT 0 99.435 0.070 100.065 ;
    RECT 0 100.135 0.070 100.765 ;
    RECT 0 100.835 0.070 101.465 ;
    RECT 0 101.535 0.070 102.165 ;
    RECT 0 102.235 0.070 102.865 ;
    RECT 0 102.935 0.070 103.565 ;
    RECT 0 103.635 0.070 104.265 ;
    RECT 0 104.335 0.070 104.965 ;
    RECT 0 105.035 0.070 105.665 ;
    RECT 0 105.735 0.070 106.365 ;
    RECT 0 106.435 0.070 107.065 ;
    RECT 0 107.135 0.070 107.765 ;
    RECT 0 107.835 0.070 108.465 ;
    RECT 0 108.535 0.070 109.165 ;
    RECT 0 109.235 0.070 109.865 ;
    RECT 0 109.935 0.070 110.565 ;
    RECT 0 110.635 0.070 111.265 ;
    RECT 0 111.335 0.070 111.965 ;
    RECT 0 112.035 0.070 112.665 ;
    RECT 0 112.735 0.070 113.365 ;
    RECT 0 113.435 0.070 114.065 ;
    RECT 0 114.135 0.070 114.765 ;
    RECT 0 114.835 0.070 115.465 ;
    RECT 0 115.535 0.070 116.165 ;
    RECT 0 116.235 0.070 116.865 ;
    RECT 0 116.935 0.070 117.565 ;
    RECT 0 117.635 0.070 118.265 ;
    RECT 0 118.335 0.070 118.965 ;
    RECT 0 119.035 0.070 119.665 ;
    RECT 0 119.735 0.070 120.365 ;
    RECT 0 120.435 0.070 121.065 ;
    RECT 0 121.135 0.070 121.765 ;
    RECT 0 121.835 0.070 122.465 ;
    RECT 0 122.535 0.070 123.165 ;
    RECT 0 123.235 0.070 123.865 ;
    RECT 0 123.935 0.070 124.565 ;
    RECT 0 124.635 0.070 125.265 ;
    RECT 0 125.335 0.070 125.965 ;
    RECT 0 126.035 0.070 126.665 ;
    RECT 0 126.735 0.070 127.365 ;
    RECT 0 127.435 0.070 128.065 ;
    RECT 0 128.135 0.070 128.765 ;
    RECT 0 128.835 0.070 129.465 ;
    RECT 0 129.535 0.070 130.165 ;
    RECT 0 130.235 0.070 130.865 ;
    RECT 0 130.935 0.070 131.565 ;
    RECT 0 131.635 0.070 132.265 ;
    RECT 0 132.335 0.070 132.965 ;
    RECT 0 133.035 0.070 133.665 ;
    RECT 0 133.735 0.070 134.365 ;
    RECT 0 134.435 0.070 135.065 ;
    RECT 0 135.135 0.070 135.765 ;
    RECT 0 135.835 0.070 136.465 ;
    RECT 0 136.535 0.070 137.165 ;
    RECT 0 137.235 0.070 137.865 ;
    RECT 0 137.935 0.070 138.565 ;
    RECT 0 138.635 0.070 139.265 ;
    RECT 0 139.335 0.070 139.965 ;
    RECT 0 140.035 0.070 140.665 ;
    RECT 0 140.735 0.070 141.365 ;
    RECT 0 141.435 0.070 142.065 ;
    RECT 0 142.135 0.070 142.765 ;
    RECT 0 142.835 0.070 143.465 ;
    RECT 0 143.535 0.070 144.165 ;
    RECT 0 144.235 0.070 144.865 ;
    RECT 0 144.935 0.070 145.565 ;
    RECT 0 145.635 0.070 146.265 ;
    RECT 0 146.335 0.070 146.965 ;
    RECT 0 147.035 0.070 147.665 ;
    RECT 0 147.735 0.070 148.365 ;
    RECT 0 148.435 0.070 149.065 ;
    RECT 0 149.135 0.070 149.765 ;
    RECT 0 149.835 0.070 150.465 ;
    RECT 0 150.535 0.070 151.165 ;
    RECT 0 151.235 0.070 151.865 ;
    RECT 0 151.935 0.070 152.565 ;
    RECT 0 152.635 0.070 153.265 ;
    RECT 0 153.335 0.070 153.965 ;
    RECT 0 154.035 0.070 154.665 ;
    RECT 0 154.735 0.070 155.365 ;
    RECT 0 155.435 0.070 156.065 ;
    RECT 0 156.135 0.070 156.765 ;
    RECT 0 156.835 0.070 157.465 ;
    RECT 0 157.535 0.070 158.165 ;
    RECT 0 158.235 0.070 158.865 ;
    RECT 0 158.935 0.070 159.565 ;
    RECT 0 159.635 0.070 160.265 ;
    RECT 0 160.335 0.070 160.965 ;
    RECT 0 161.035 0.070 161.665 ;
    RECT 0 161.735 0.070 162.365 ;
    RECT 0 162.435 0.070 163.065 ;
    RECT 0 163.135 0.070 163.765 ;
    RECT 0 163.835 0.070 164.465 ;
    RECT 0 164.535 0.070 165.165 ;
    RECT 0 165.235 0.070 165.865 ;
    RECT 0 165.935 0.070 166.565 ;
    RECT 0 166.635 0.070 167.265 ;
    RECT 0 167.335 0.070 167.965 ;
    RECT 0 168.035 0.070 168.665 ;
    RECT 0 168.735 0.070 169.365 ;
    RECT 0 169.435 0.070 170.065 ;
    RECT 0 170.135 0.070 170.765 ;
    RECT 0 170.835 0.070 171.465 ;
    RECT 0 171.535 0.070 172.165 ;
    RECT 0 172.235 0.070 172.865 ;
    RECT 0 172.935 0.070 173.565 ;
    RECT 0 173.635 0.070 174.265 ;
    RECT 0 174.335 0.070 174.965 ;
    RECT 0 175.035 0.070 175.665 ;
    RECT 0 175.735 0.070 176.365 ;
    RECT 0 176.435 0.070 177.065 ;
    RECT 0 177.135 0.070 177.765 ;
    RECT 0 177.835 0.070 178.465 ;
    RECT 0 178.535 0.070 179.165 ;
    RECT 0 179.235 0.070 179.865 ;
    RECT 0 179.935 0.070 180.565 ;
    RECT 0 180.635 0.070 181.265 ;
    RECT 0 181.335 0.070 181.965 ;
    RECT 0 182.035 0.070 182.665 ;
    RECT 0 182.735 0.070 183.365 ;
    RECT 0 183.435 0.070 184.065 ;
    RECT 0 184.135 0.070 184.765 ;
    RECT 0 184.835 0.070 185.465 ;
    RECT 0 185.535 0.070 186.165 ;
    RECT 0 186.235 0.070 186.865 ;
    RECT 0 186.935 0.070 187.565 ;
    RECT 0 187.635 0.070 188.265 ;
    RECT 0 188.335 0.070 188.965 ;
    RECT 0 189.035 0.070 189.665 ;
    RECT 0 189.735 0.070 190.365 ;
    RECT 0 190.435 0.070 191.065 ;
    RECT 0 191.135 0.070 191.765 ;
    RECT 0 191.835 0.070 192.465 ;
    RECT 0 192.535 0.070 193.165 ;
    RECT 0 193.235 0.070 193.865 ;
    RECT 0 193.935 0.070 194.565 ;
    RECT 0 194.635 0.070 195.265 ;
    RECT 0 195.335 0.070 195.965 ;
    RECT 0 196.035 0.070 196.665 ;
    RECT 0 196.735 0.070 197.365 ;
    RECT 0 197.435 0.070 198.065 ;
    RECT 0 198.135 0.070 198.765 ;
    RECT 0 198.835 0.070 199.465 ;
    RECT 0 199.535 0.070 200.165 ;
    RECT 0 200.235 0.070 200.865 ;
    RECT 0 200.935 0.070 201.565 ;
    RECT 0 201.635 0.070 202.265 ;
    RECT 0 202.335 0.070 202.965 ;
    RECT 0 203.035 0.070 203.665 ;
    RECT 0 203.735 0.070 204.365 ;
    RECT 0 204.435 0.070 205.065 ;
    RECT 0 205.135 0.070 205.765 ;
    RECT 0 205.835 0.070 206.465 ;
    RECT 0 206.535 0.070 207.165 ;
    RECT 0 207.235 0.070 207.865 ;
    RECT 0 207.935 0.070 208.565 ;
    RECT 0 208.635 0.070 209.265 ;
    RECT 0 209.335 0.070 209.965 ;
    RECT 0 210.035 0.070 210.665 ;
    RECT 0 210.735 0.070 211.365 ;
    RECT 0 211.435 0.070 212.065 ;
    RECT 0 212.135 0.070 212.765 ;
    RECT 0 212.835 0.070 213.465 ;
    RECT 0 213.535 0.070 214.165 ;
    RECT 0 214.235 0.070 214.865 ;
    RECT 0 214.935 0.070 215.565 ;
    RECT 0 215.635 0.070 216.265 ;
    RECT 0 216.335 0.070 216.965 ;
    RECT 0 217.035 0.070 217.665 ;
    RECT 0 217.735 0.070 218.365 ;
    RECT 0 218.435 0.070 219.065 ;
    RECT 0 219.135 0.070 219.765 ;
    RECT 0 219.835 0.070 220.465 ;
    RECT 0 220.535 0.070 221.165 ;
    RECT 0 221.235 0.070 221.865 ;
    RECT 0 221.935 0.070 222.565 ;
    RECT 0 222.635 0.070 223.265 ;
    RECT 0 223.335 0.070 223.965 ;
    RECT 0 224.035 0.070 224.665 ;
    RECT 0 224.735 0.070 225.365 ;
    RECT 0 225.435 0.070 226.065 ;
    RECT 0 226.135 0.070 226.765 ;
    RECT 0 226.835 0.070 227.465 ;
    RECT 0 227.535 0.070 228.165 ;
    RECT 0 228.235 0.070 228.865 ;
    RECT 0 228.935 0.070 229.565 ;
    RECT 0 229.635 0.070 230.265 ;
    RECT 0 230.335 0.070 230.965 ;
    RECT 0 231.035 0.070 231.665 ;
    RECT 0 231.735 0.070 232.365 ;
    RECT 0 232.435 0.070 233.065 ;
    RECT 0 233.135 0.070 233.765 ;
    RECT 0 233.835 0.070 234.465 ;
    RECT 0 234.535 0.070 235.165 ;
    RECT 0 235.235 0.070 235.865 ;
    RECT 0 235.935 0.070 236.565 ;
    RECT 0 236.635 0.070 237.265 ;
    RECT 0 237.335 0.070 237.965 ;
    RECT 0 238.035 0.070 238.665 ;
    RECT 0 238.735 0.070 239.365 ;
    RECT 0 239.435 0.070 240.065 ;
    RECT 0 240.135 0.070 240.765 ;
    RECT 0 240.835 0.070 241.465 ;
    RECT 0 241.535 0.070 242.165 ;
    RECT 0 242.235 0.070 242.865 ;
    RECT 0 242.935 0.070 243.565 ;
    RECT 0 243.635 0.070 244.265 ;
    RECT 0 244.335 0.070 244.965 ;
    RECT 0 245.035 0.070 245.665 ;
    RECT 0 245.735 0.070 246.365 ;
    RECT 0 246.435 0.070 247.065 ;
    RECT 0 247.135 0.070 247.765 ;
    RECT 0 247.835 0.070 248.465 ;
    RECT 0 248.535 0.070 249.165 ;
    RECT 0 249.235 0.070 249.865 ;
    RECT 0 249.935 0.070 250.565 ;
    RECT 0 250.635 0.070 251.265 ;
    RECT 0 251.335 0.070 251.965 ;
    RECT 0 252.035 0.070 252.665 ;
    RECT 0 252.735 0.070 253.365 ;
    RECT 0 253.435 0.070 254.065 ;
    RECT 0 254.135 0.070 254.765 ;
    RECT 0 254.835 0.070 255.465 ;
    RECT 0 255.535 0.070 256.165 ;
    RECT 0 256.235 0.070 256.865 ;
    RECT 0 256.935 0.070 257.565 ;
    RECT 0 257.635 0.070 258.265 ;
    RECT 0 258.335 0.070 258.965 ;
    RECT 0 259.035 0.070 259.665 ;
    RECT 0 259.735 0.070 260.365 ;
    RECT 0 260.435 0.070 261.065 ;
    RECT 0 261.135 0.070 261.765 ;
    RECT 0 261.835 0.070 262.465 ;
    RECT 0 262.535 0.070 263.165 ;
    RECT 0 263.235 0.070 263.865 ;
    RECT 0 263.935 0.070 264.565 ;
    RECT 0 264.635 0.070 265.265 ;
    RECT 0 265.335 0.070 265.965 ;
    RECT 0 266.035 0.070 266.665 ;
    RECT 0 266.735 0.070 267.365 ;
    RECT 0 267.435 0.070 268.065 ;
    RECT 0 268.135 0.070 268.765 ;
    RECT 0 268.835 0.070 269.465 ;
    RECT 0 269.535 0.070 270.165 ;
    RECT 0 270.235 0.070 270.865 ;
    RECT 0 270.935 0.070 271.565 ;
    RECT 0 271.635 0.070 272.265 ;
    RECT 0 272.335 0.070 272.965 ;
    RECT 0 273.035 0.070 273.665 ;
    RECT 0 273.735 0.070 274.365 ;
    RECT 0 274.435 0.070 275.065 ;
    RECT 0 275.135 0.070 275.765 ;
    RECT 0 275.835 0.070 276.465 ;
    RECT 0 276.535 0.070 277.165 ;
    RECT 0 277.235 0.070 277.865 ;
    RECT 0 277.935 0.070 278.565 ;
    RECT 0 278.635 0.070 279.265 ;
    RECT 0 279.335 0.070 279.965 ;
    RECT 0 280.035 0.070 280.665 ;
    RECT 0 280.735 0.070 281.365 ;
    RECT 0 281.435 0.070 282.065 ;
    RECT 0 282.135 0.070 282.765 ;
    RECT 0 282.835 0.070 283.465 ;
    RECT 0 283.535 0.070 284.165 ;
    RECT 0 284.235 0.070 284.865 ;
    RECT 0 284.935 0.070 285.565 ;
    RECT 0 285.635 0.070 286.265 ;
    RECT 0 286.335 0.070 286.965 ;
    RECT 0 287.035 0.070 287.665 ;
    RECT 0 287.735 0.070 288.365 ;
    RECT 0 288.435 0.070 289.065 ;
    RECT 0 289.135 0.070 289.765 ;
    RECT 0 289.835 0.070 290.465 ;
    RECT 0 290.535 0.070 291.165 ;
    RECT 0 291.235 0.070 291.865 ;
    RECT 0 291.935 0.070 292.565 ;
    RECT 0 292.635 0.070 293.265 ;
    RECT 0 293.335 0.070 293.965 ;
    RECT 0 294.035 0.070 294.665 ;
    RECT 0 294.735 0.070 295.365 ;
    RECT 0 295.435 0.070 296.065 ;
    RECT 0 296.135 0.070 296.765 ;
    RECT 0 296.835 0.070 297.465 ;
    RECT 0 297.535 0.070 298.165 ;
    RECT 0 298.235 0.070 298.865 ;
    RECT 0 298.935 0.070 299.565 ;
    RECT 0 299.635 0.070 300.265 ;
    RECT 0 300.335 0.070 300.965 ;
    RECT 0 301.035 0.070 301.665 ;
    RECT 0 301.735 0.070 302.365 ;
    RECT 0 302.435 0.070 303.065 ;
    RECT 0 303.135 0.070 303.765 ;
    RECT 0 303.835 0.070 304.465 ;
    RECT 0 304.535 0.070 305.165 ;
    RECT 0 305.235 0.070 305.865 ;
    RECT 0 305.935 0.070 306.565 ;
    RECT 0 306.635 0.070 307.265 ;
    RECT 0 307.335 0.070 307.965 ;
    RECT 0 308.035 0.070 308.665 ;
    RECT 0 308.735 0.070 309.365 ;
    RECT 0 309.435 0.070 310.065 ;
    RECT 0 310.135 0.070 310.765 ;
    RECT 0 310.835 0.070 311.465 ;
    RECT 0 311.535 0.070 312.165 ;
    RECT 0 312.235 0.070 312.865 ;
    RECT 0 312.935 0.070 313.565 ;
    RECT 0 313.635 0.070 314.265 ;
    RECT 0 314.335 0.070 314.965 ;
    RECT 0 315.035 0.070 315.665 ;
    RECT 0 315.735 0.070 316.365 ;
    RECT 0 316.435 0.070 317.065 ;
    RECT 0 317.135 0.070 317.765 ;
    RECT 0 317.835 0.070 318.465 ;
    RECT 0 318.535 0.070 319.165 ;
    RECT 0 319.235 0.070 319.865 ;
    RECT 0 319.935 0.070 320.565 ;
    RECT 0 320.635 0.070 321.265 ;
    RECT 0 321.335 0.070 321.965 ;
    RECT 0 322.035 0.070 322.665 ;
    RECT 0 322.735 0.070 323.365 ;
    RECT 0 323.435 0.070 324.065 ;
    RECT 0 324.135 0.070 324.765 ;
    RECT 0 324.835 0.070 325.465 ;
    RECT 0 325.535 0.070 326.165 ;
    RECT 0 326.235 0.070 326.865 ;
    RECT 0 326.935 0.070 327.565 ;
    RECT 0 327.635 0.070 328.265 ;
    RECT 0 328.335 0.070 328.965 ;
    RECT 0 329.035 0.070 329.665 ;
    RECT 0 329.735 0.070 330.365 ;
    RECT 0 330.435 0.070 331.065 ;
    RECT 0 331.135 0.070 331.765 ;
    RECT 0 331.835 0.070 332.465 ;
    RECT 0 332.535 0.070 333.165 ;
    RECT 0 333.235 0.070 333.865 ;
    RECT 0 333.935 0.070 334.565 ;
    RECT 0 334.635 0.070 335.265 ;
    RECT 0 335.335 0.070 335.965 ;
    RECT 0 336.035 0.070 336.665 ;
    RECT 0 336.735 0.070 337.365 ;
    RECT 0 337.435 0.070 338.065 ;
    RECT 0 338.135 0.070 338.765 ;
    RECT 0 338.835 0.070 339.465 ;
    RECT 0 339.535 0.070 340.165 ;
    RECT 0 340.235 0.070 340.865 ;
    RECT 0 340.935 0.070 341.565 ;
    RECT 0 341.635 0.070 342.265 ;
    RECT 0 342.335 0.070 342.965 ;
    RECT 0 343.035 0.070 343.665 ;
    RECT 0 343.735 0.070 344.365 ;
    RECT 0 344.435 0.070 345.065 ;
    RECT 0 345.135 0.070 345.765 ;
    RECT 0 345.835 0.070 346.465 ;
    RECT 0 346.535 0.070 347.165 ;
    RECT 0 347.235 0.070 347.865 ;
    RECT 0 347.935 0.070 348.565 ;
    RECT 0 348.635 0.070 349.265 ;
    RECT 0 349.335 0.070 349.965 ;
    RECT 0 350.035 0.070 350.665 ;
    RECT 0 350.735 0.070 351.365 ;
    RECT 0 351.435 0.070 352.065 ;
    RECT 0 352.135 0.070 352.765 ;
    RECT 0 352.835 0.070 353.465 ;
    RECT 0 353.535 0.070 354.165 ;
    RECT 0 354.235 0.070 354.865 ;
    RECT 0 354.935 0.070 355.565 ;
    RECT 0 355.635 0.070 356.265 ;
    RECT 0 356.335 0.070 356.965 ;
    RECT 0 357.035 0.070 357.665 ;
    RECT 0 357.735 0.070 358.365 ;
    RECT 0 358.435 0.070 359.065 ;
    RECT 0 359.135 0.070 407.085 ;
    RECT 0 407.155 0.070 407.785 ;
    RECT 0 407.855 0.070 408.485 ;
    RECT 0 408.555 0.070 409.185 ;
    RECT 0 409.255 0.070 409.885 ;
    RECT 0 409.955 0.070 410.585 ;
    RECT 0 410.655 0.070 411.285 ;
    RECT 0 411.355 0.070 411.985 ;
    RECT 0 412.055 0.070 412.685 ;
    RECT 0 412.755 0.070 413.385 ;
    RECT 0 413.455 0.070 414.085 ;
    RECT 0 414.155 0.070 414.785 ;
    RECT 0 414.855 0.070 415.485 ;
    RECT 0 415.555 0.070 416.185 ;
    RECT 0 416.255 0.070 416.885 ;
    RECT 0 416.955 0.070 417.585 ;
    RECT 0 417.655 0.070 418.285 ;
    RECT 0 418.355 0.070 418.985 ;
    RECT 0 419.055 0.070 419.685 ;
    RECT 0 419.755 0.070 420.385 ;
    RECT 0 420.455 0.070 421.085 ;
    RECT 0 421.155 0.070 421.785 ;
    RECT 0 421.855 0.070 422.485 ;
    RECT 0 422.555 0.070 423.185 ;
    RECT 0 423.255 0.070 423.885 ;
    RECT 0 423.955 0.070 424.585 ;
    RECT 0 424.655 0.070 425.285 ;
    RECT 0 425.355 0.070 425.985 ;
    RECT 0 426.055 0.070 426.685 ;
    RECT 0 426.755 0.070 427.385 ;
    RECT 0 427.455 0.070 428.085 ;
    RECT 0 428.155 0.070 428.785 ;
    RECT 0 428.855 0.070 429.485 ;
    RECT 0 429.555 0.070 430.185 ;
    RECT 0 430.255 0.070 430.885 ;
    RECT 0 430.955 0.070 431.585 ;
    RECT 0 431.655 0.070 432.285 ;
    RECT 0 432.355 0.070 432.985 ;
    RECT 0 433.055 0.070 433.685 ;
    RECT 0 433.755 0.070 434.385 ;
    RECT 0 434.455 0.070 435.085 ;
    RECT 0 435.155 0.070 435.785 ;
    RECT 0 435.855 0.070 436.485 ;
    RECT 0 436.555 0.070 437.185 ;
    RECT 0 437.255 0.070 437.885 ;
    RECT 0 437.955 0.070 438.585 ;
    RECT 0 438.655 0.070 439.285 ;
    RECT 0 439.355 0.070 439.985 ;
    RECT 0 440.055 0.070 440.685 ;
    RECT 0 440.755 0.070 441.385 ;
    RECT 0 441.455 0.070 442.085 ;
    RECT 0 442.155 0.070 442.785 ;
    RECT 0 442.855 0.070 443.485 ;
    RECT 0 443.555 0.070 444.185 ;
    RECT 0 444.255 0.070 444.885 ;
    RECT 0 444.955 0.070 445.585 ;
    RECT 0 445.655 0.070 446.285 ;
    RECT 0 446.355 0.070 446.985 ;
    RECT 0 447.055 0.070 447.685 ;
    RECT 0 447.755 0.070 448.385 ;
    RECT 0 448.455 0.070 449.085 ;
    RECT 0 449.155 0.070 449.785 ;
    RECT 0 449.855 0.070 450.485 ;
    RECT 0 450.555 0.070 451.185 ;
    RECT 0 451.255 0.070 451.885 ;
    RECT 0 451.955 0.070 452.585 ;
    RECT 0 452.655 0.070 453.285 ;
    RECT 0 453.355 0.070 453.985 ;
    RECT 0 454.055 0.070 454.685 ;
    RECT 0 454.755 0.070 455.385 ;
    RECT 0 455.455 0.070 456.085 ;
    RECT 0 456.155 0.070 456.785 ;
    RECT 0 456.855 0.070 457.485 ;
    RECT 0 457.555 0.070 458.185 ;
    RECT 0 458.255 0.070 458.885 ;
    RECT 0 458.955 0.070 459.585 ;
    RECT 0 459.655 0.070 460.285 ;
    RECT 0 460.355 0.070 460.985 ;
    RECT 0 461.055 0.070 461.685 ;
    RECT 0 461.755 0.070 462.385 ;
    RECT 0 462.455 0.070 463.085 ;
    RECT 0 463.155 0.070 463.785 ;
    RECT 0 463.855 0.070 464.485 ;
    RECT 0 464.555 0.070 465.185 ;
    RECT 0 465.255 0.070 465.885 ;
    RECT 0 465.955 0.070 466.585 ;
    RECT 0 466.655 0.070 467.285 ;
    RECT 0 467.355 0.070 467.985 ;
    RECT 0 468.055 0.070 468.685 ;
    RECT 0 468.755 0.070 469.385 ;
    RECT 0 469.455 0.070 470.085 ;
    RECT 0 470.155 0.070 470.785 ;
    RECT 0 470.855 0.070 471.485 ;
    RECT 0 471.555 0.070 472.185 ;
    RECT 0 472.255 0.070 472.885 ;
    RECT 0 472.955 0.070 473.585 ;
    RECT 0 473.655 0.070 474.285 ;
    RECT 0 474.355 0.070 474.985 ;
    RECT 0 475.055 0.070 475.685 ;
    RECT 0 475.755 0.070 476.385 ;
    RECT 0 476.455 0.070 477.085 ;
    RECT 0 477.155 0.070 477.785 ;
    RECT 0 477.855 0.070 478.485 ;
    RECT 0 478.555 0.070 479.185 ;
    RECT 0 479.255 0.070 479.885 ;
    RECT 0 479.955 0.070 480.585 ;
    RECT 0 480.655 0.070 481.285 ;
    RECT 0 481.355 0.070 481.985 ;
    RECT 0 482.055 0.070 482.685 ;
    RECT 0 482.755 0.070 483.385 ;
    RECT 0 483.455 0.070 484.085 ;
    RECT 0 484.155 0.070 484.785 ;
    RECT 0 484.855 0.070 485.485 ;
    RECT 0 485.555 0.070 486.185 ;
    RECT 0 486.255 0.070 486.885 ;
    RECT 0 486.955 0.070 487.585 ;
    RECT 0 487.655 0.070 488.285 ;
    RECT 0 488.355 0.070 488.985 ;
    RECT 0 489.055 0.070 489.685 ;
    RECT 0 489.755 0.070 490.385 ;
    RECT 0 490.455 0.070 491.085 ;
    RECT 0 491.155 0.070 491.785 ;
    RECT 0 491.855 0.070 492.485 ;
    RECT 0 492.555 0.070 493.185 ;
    RECT 0 493.255 0.070 493.885 ;
    RECT 0 493.955 0.070 494.585 ;
    RECT 0 494.655 0.070 495.285 ;
    RECT 0 495.355 0.070 495.985 ;
    RECT 0 496.055 0.070 496.685 ;
    RECT 0 496.755 0.070 497.385 ;
    RECT 0 497.455 0.070 498.085 ;
    RECT 0 498.155 0.070 498.785 ;
    RECT 0 498.855 0.070 499.485 ;
    RECT 0 499.555 0.070 500.185 ;
    RECT 0 500.255 0.070 500.885 ;
    RECT 0 500.955 0.070 501.585 ;
    RECT 0 501.655 0.070 502.285 ;
    RECT 0 502.355 0.070 502.985 ;
    RECT 0 503.055 0.070 503.685 ;
    RECT 0 503.755 0.070 504.385 ;
    RECT 0 504.455 0.070 505.085 ;
    RECT 0 505.155 0.070 505.785 ;
    RECT 0 505.855 0.070 506.485 ;
    RECT 0 506.555 0.070 507.185 ;
    RECT 0 507.255 0.070 507.885 ;
    RECT 0 507.955 0.070 508.585 ;
    RECT 0 508.655 0.070 509.285 ;
    RECT 0 509.355 0.070 509.985 ;
    RECT 0 510.055 0.070 510.685 ;
    RECT 0 510.755 0.070 511.385 ;
    RECT 0 511.455 0.070 512.085 ;
    RECT 0 512.155 0.070 512.785 ;
    RECT 0 512.855 0.070 513.485 ;
    RECT 0 513.555 0.070 514.185 ;
    RECT 0 514.255 0.070 514.885 ;
    RECT 0 514.955 0.070 515.585 ;
    RECT 0 515.655 0.070 516.285 ;
    RECT 0 516.355 0.070 516.985 ;
    RECT 0 517.055 0.070 517.685 ;
    RECT 0 517.755 0.070 518.385 ;
    RECT 0 518.455 0.070 519.085 ;
    RECT 0 519.155 0.070 519.785 ;
    RECT 0 519.855 0.070 520.485 ;
    RECT 0 520.555 0.070 521.185 ;
    RECT 0 521.255 0.070 521.885 ;
    RECT 0 521.955 0.070 522.585 ;
    RECT 0 522.655 0.070 523.285 ;
    RECT 0 523.355 0.070 523.985 ;
    RECT 0 524.055 0.070 524.685 ;
    RECT 0 524.755 0.070 525.385 ;
    RECT 0 525.455 0.070 526.085 ;
    RECT 0 526.155 0.070 526.785 ;
    RECT 0 526.855 0.070 527.485 ;
    RECT 0 527.555 0.070 528.185 ;
    RECT 0 528.255 0.070 528.885 ;
    RECT 0 528.955 0.070 529.585 ;
    RECT 0 529.655 0.070 530.285 ;
    RECT 0 530.355 0.070 530.985 ;
    RECT 0 531.055 0.070 531.685 ;
    RECT 0 531.755 0.070 532.385 ;
    RECT 0 532.455 0.070 533.085 ;
    RECT 0 533.155 0.070 533.785 ;
    RECT 0 533.855 0.070 534.485 ;
    RECT 0 534.555 0.070 535.185 ;
    RECT 0 535.255 0.070 535.885 ;
    RECT 0 535.955 0.070 536.585 ;
    RECT 0 536.655 0.070 537.285 ;
    RECT 0 537.355 0.070 537.985 ;
    RECT 0 538.055 0.070 538.685 ;
    RECT 0 538.755 0.070 539.385 ;
    RECT 0 539.455 0.070 540.085 ;
    RECT 0 540.155 0.070 540.785 ;
    RECT 0 540.855 0.070 541.485 ;
    RECT 0 541.555 0.070 542.185 ;
    RECT 0 542.255 0.070 542.885 ;
    RECT 0 542.955 0.070 543.585 ;
    RECT 0 543.655 0.070 544.285 ;
    RECT 0 544.355 0.070 544.985 ;
    RECT 0 545.055 0.070 545.685 ;
    RECT 0 545.755 0.070 546.385 ;
    RECT 0 546.455 0.070 547.085 ;
    RECT 0 547.155 0.070 547.785 ;
    RECT 0 547.855 0.070 548.485 ;
    RECT 0 548.555 0.070 549.185 ;
    RECT 0 549.255 0.070 549.885 ;
    RECT 0 549.955 0.070 550.585 ;
    RECT 0 550.655 0.070 551.285 ;
    RECT 0 551.355 0.070 551.985 ;
    RECT 0 552.055 0.070 552.685 ;
    RECT 0 552.755 0.070 553.385 ;
    RECT 0 553.455 0.070 554.085 ;
    RECT 0 554.155 0.070 554.785 ;
    RECT 0 554.855 0.070 555.485 ;
    RECT 0 555.555 0.070 556.185 ;
    RECT 0 556.255 0.070 556.885 ;
    RECT 0 556.955 0.070 557.585 ;
    RECT 0 557.655 0.070 558.285 ;
    RECT 0 558.355 0.070 558.985 ;
    RECT 0 559.055 0.070 559.685 ;
    RECT 0 559.755 0.070 560.385 ;
    RECT 0 560.455 0.070 561.085 ;
    RECT 0 561.155 0.070 561.785 ;
    RECT 0 561.855 0.070 562.485 ;
    RECT 0 562.555 0.070 563.185 ;
    RECT 0 563.255 0.070 563.885 ;
    RECT 0 563.955 0.070 564.585 ;
    RECT 0 564.655 0.070 565.285 ;
    RECT 0 565.355 0.070 565.985 ;
    RECT 0 566.055 0.070 566.685 ;
    RECT 0 566.755 0.070 567.385 ;
    RECT 0 567.455 0.070 568.085 ;
    RECT 0 568.155 0.070 568.785 ;
    RECT 0 568.855 0.070 569.485 ;
    RECT 0 569.555 0.070 570.185 ;
    RECT 0 570.255 0.070 570.885 ;
    RECT 0 570.955 0.070 571.585 ;
    RECT 0 571.655 0.070 572.285 ;
    RECT 0 572.355 0.070 572.985 ;
    RECT 0 573.055 0.070 573.685 ;
    RECT 0 573.755 0.070 574.385 ;
    RECT 0 574.455 0.070 575.085 ;
    RECT 0 575.155 0.070 575.785 ;
    RECT 0 575.855 0.070 576.485 ;
    RECT 0 576.555 0.070 577.185 ;
    RECT 0 577.255 0.070 577.885 ;
    RECT 0 577.955 0.070 578.585 ;
    RECT 0 578.655 0.070 579.285 ;
    RECT 0 579.355 0.070 579.985 ;
    RECT 0 580.055 0.070 580.685 ;
    RECT 0 580.755 0.070 581.385 ;
    RECT 0 581.455 0.070 582.085 ;
    RECT 0 582.155 0.070 582.785 ;
    RECT 0 582.855 0.070 583.485 ;
    RECT 0 583.555 0.070 584.185 ;
    RECT 0 584.255 0.070 584.885 ;
    RECT 0 584.955 0.070 585.585 ;
    RECT 0 585.655 0.070 586.285 ;
    RECT 0 586.355 0.070 586.985 ;
    RECT 0 587.055 0.070 587.685 ;
    RECT 0 587.755 0.070 588.385 ;
    RECT 0 588.455 0.070 589.085 ;
    RECT 0 589.155 0.070 589.785 ;
    RECT 0 589.855 0.070 590.485 ;
    RECT 0 590.555 0.070 591.185 ;
    RECT 0 591.255 0.070 591.885 ;
    RECT 0 591.955 0.070 592.585 ;
    RECT 0 592.655 0.070 593.285 ;
    RECT 0 593.355 0.070 593.985 ;
    RECT 0 594.055 0.070 594.685 ;
    RECT 0 594.755 0.070 595.385 ;
    RECT 0 595.455 0.070 596.085 ;
    RECT 0 596.155 0.070 596.785 ;
    RECT 0 596.855 0.070 597.485 ;
    RECT 0 597.555 0.070 598.185 ;
    RECT 0 598.255 0.070 598.885 ;
    RECT 0 598.955 0.070 599.585 ;
    RECT 0 599.655 0.070 600.285 ;
    RECT 0 600.355 0.070 600.985 ;
    RECT 0 601.055 0.070 601.685 ;
    RECT 0 601.755 0.070 602.385 ;
    RECT 0 602.455 0.070 603.085 ;
    RECT 0 603.155 0.070 603.785 ;
    RECT 0 603.855 0.070 604.485 ;
    RECT 0 604.555 0.070 605.185 ;
    RECT 0 605.255 0.070 605.885 ;
    RECT 0 605.955 0.070 606.585 ;
    RECT 0 606.655 0.070 607.285 ;
    RECT 0 607.355 0.070 607.985 ;
    RECT 0 608.055 0.070 608.685 ;
    RECT 0 608.755 0.070 609.385 ;
    RECT 0 609.455 0.070 610.085 ;
    RECT 0 610.155 0.070 610.785 ;
    RECT 0 610.855 0.070 611.485 ;
    RECT 0 611.555 0.070 612.185 ;
    RECT 0 612.255 0.070 612.885 ;
    RECT 0 612.955 0.070 613.585 ;
    RECT 0 613.655 0.070 614.285 ;
    RECT 0 614.355 0.070 614.985 ;
    RECT 0 615.055 0.070 615.685 ;
    RECT 0 615.755 0.070 616.385 ;
    RECT 0 616.455 0.070 617.085 ;
    RECT 0 617.155 0.070 617.785 ;
    RECT 0 617.855 0.070 618.485 ;
    RECT 0 618.555 0.070 619.185 ;
    RECT 0 619.255 0.070 619.885 ;
    RECT 0 619.955 0.070 620.585 ;
    RECT 0 620.655 0.070 621.285 ;
    RECT 0 621.355 0.070 621.985 ;
    RECT 0 622.055 0.070 622.685 ;
    RECT 0 622.755 0.070 623.385 ;
    RECT 0 623.455 0.070 624.085 ;
    RECT 0 624.155 0.070 624.785 ;
    RECT 0 624.855 0.070 625.485 ;
    RECT 0 625.555 0.070 626.185 ;
    RECT 0 626.255 0.070 626.885 ;
    RECT 0 626.955 0.070 627.585 ;
    RECT 0 627.655 0.070 628.285 ;
    RECT 0 628.355 0.070 628.985 ;
    RECT 0 629.055 0.070 629.685 ;
    RECT 0 629.755 0.070 630.385 ;
    RECT 0 630.455 0.070 631.085 ;
    RECT 0 631.155 0.070 631.785 ;
    RECT 0 631.855 0.070 632.485 ;
    RECT 0 632.555 0.070 633.185 ;
    RECT 0 633.255 0.070 633.885 ;
    RECT 0 633.955 0.070 634.585 ;
    RECT 0 634.655 0.070 635.285 ;
    RECT 0 635.355 0.070 635.985 ;
    RECT 0 636.055 0.070 636.685 ;
    RECT 0 636.755 0.070 637.385 ;
    RECT 0 637.455 0.070 638.085 ;
    RECT 0 638.155 0.070 638.785 ;
    RECT 0 638.855 0.070 639.485 ;
    RECT 0 639.555 0.070 640.185 ;
    RECT 0 640.255 0.070 640.885 ;
    RECT 0 640.955 0.070 641.585 ;
    RECT 0 641.655 0.070 642.285 ;
    RECT 0 642.355 0.070 642.985 ;
    RECT 0 643.055 0.070 643.685 ;
    RECT 0 643.755 0.070 644.385 ;
    RECT 0 644.455 0.070 645.085 ;
    RECT 0 645.155 0.070 645.785 ;
    RECT 0 645.855 0.070 646.485 ;
    RECT 0 646.555 0.070 647.185 ;
    RECT 0 647.255 0.070 647.885 ;
    RECT 0 647.955 0.070 648.585 ;
    RECT 0 648.655 0.070 649.285 ;
    RECT 0 649.355 0.070 649.985 ;
    RECT 0 650.055 0.070 650.685 ;
    RECT 0 650.755 0.070 651.385 ;
    RECT 0 651.455 0.070 652.085 ;
    RECT 0 652.155 0.070 652.785 ;
    RECT 0 652.855 0.070 653.485 ;
    RECT 0 653.555 0.070 654.185 ;
    RECT 0 654.255 0.070 654.885 ;
    RECT 0 654.955 0.070 655.585 ;
    RECT 0 655.655 0.070 656.285 ;
    RECT 0 656.355 0.070 656.985 ;
    RECT 0 657.055 0.070 657.685 ;
    RECT 0 657.755 0.070 658.385 ;
    RECT 0 658.455 0.070 659.085 ;
    RECT 0 659.155 0.070 659.785 ;
    RECT 0 659.855 0.070 660.485 ;
    RECT 0 660.555 0.070 661.185 ;
    RECT 0 661.255 0.070 661.885 ;
    RECT 0 661.955 0.070 662.585 ;
    RECT 0 662.655 0.070 663.285 ;
    RECT 0 663.355 0.070 663.985 ;
    RECT 0 664.055 0.070 664.685 ;
    RECT 0 664.755 0.070 665.385 ;
    RECT 0 665.455 0.070 666.085 ;
    RECT 0 666.155 0.070 666.785 ;
    RECT 0 666.855 0.070 667.485 ;
    RECT 0 667.555 0.070 668.185 ;
    RECT 0 668.255 0.070 668.885 ;
    RECT 0 668.955 0.070 669.585 ;
    RECT 0 669.655 0.070 670.285 ;
    RECT 0 670.355 0.070 670.985 ;
    RECT 0 671.055 0.070 671.685 ;
    RECT 0 671.755 0.070 672.385 ;
    RECT 0 672.455 0.070 673.085 ;
    RECT 0 673.155 0.070 673.785 ;
    RECT 0 673.855 0.070 674.485 ;
    RECT 0 674.555 0.070 675.185 ;
    RECT 0 675.255 0.070 675.885 ;
    RECT 0 675.955 0.070 676.585 ;
    RECT 0 676.655 0.070 677.285 ;
    RECT 0 677.355 0.070 677.985 ;
    RECT 0 678.055 0.070 678.685 ;
    RECT 0 678.755 0.070 679.385 ;
    RECT 0 679.455 0.070 680.085 ;
    RECT 0 680.155 0.070 680.785 ;
    RECT 0 680.855 0.070 681.485 ;
    RECT 0 681.555 0.070 682.185 ;
    RECT 0 682.255 0.070 682.885 ;
    RECT 0 682.955 0.070 683.585 ;
    RECT 0 683.655 0.070 684.285 ;
    RECT 0 684.355 0.070 684.985 ;
    RECT 0 685.055 0.070 685.685 ;
    RECT 0 685.755 0.070 686.385 ;
    RECT 0 686.455 0.070 687.085 ;
    RECT 0 687.155 0.070 687.785 ;
    RECT 0 687.855 0.070 688.485 ;
    RECT 0 688.555 0.070 689.185 ;
    RECT 0 689.255 0.070 689.885 ;
    RECT 0 689.955 0.070 690.585 ;
    RECT 0 690.655 0.070 691.285 ;
    RECT 0 691.355 0.070 691.985 ;
    RECT 0 692.055 0.070 692.685 ;
    RECT 0 692.755 0.070 693.385 ;
    RECT 0 693.455 0.070 694.085 ;
    RECT 0 694.155 0.070 694.785 ;
    RECT 0 694.855 0.070 695.485 ;
    RECT 0 695.555 0.070 696.185 ;
    RECT 0 696.255 0.070 696.885 ;
    RECT 0 696.955 0.070 697.585 ;
    RECT 0 697.655 0.070 698.285 ;
    RECT 0 698.355 0.070 698.985 ;
    RECT 0 699.055 0.070 699.685 ;
    RECT 0 699.755 0.070 700.385 ;
    RECT 0 700.455 0.070 701.085 ;
    RECT 0 701.155 0.070 701.785 ;
    RECT 0 701.855 0.070 702.485 ;
    RECT 0 702.555 0.070 703.185 ;
    RECT 0 703.255 0.070 703.885 ;
    RECT 0 703.955 0.070 704.585 ;
    RECT 0 704.655 0.070 705.285 ;
    RECT 0 705.355 0.070 705.985 ;
    RECT 0 706.055 0.070 706.685 ;
    RECT 0 706.755 0.070 707.385 ;
    RECT 0 707.455 0.070 708.085 ;
    RECT 0 708.155 0.070 708.785 ;
    RECT 0 708.855 0.070 709.485 ;
    RECT 0 709.555 0.070 710.185 ;
    RECT 0 710.255 0.070 710.885 ;
    RECT 0 710.955 0.070 711.585 ;
    RECT 0 711.655 0.070 712.285 ;
    RECT 0 712.355 0.070 712.985 ;
    RECT 0 713.055 0.070 713.685 ;
    RECT 0 713.755 0.070 714.385 ;
    RECT 0 714.455 0.070 715.085 ;
    RECT 0 715.155 0.070 715.785 ;
    RECT 0 715.855 0.070 716.485 ;
    RECT 0 716.555 0.070 717.185 ;
    RECT 0 717.255 0.070 717.885 ;
    RECT 0 717.955 0.070 718.585 ;
    RECT 0 718.655 0.070 719.285 ;
    RECT 0 719.355 0.070 719.985 ;
    RECT 0 720.055 0.070 720.685 ;
    RECT 0 720.755 0.070 721.385 ;
    RECT 0 721.455 0.070 722.085 ;
    RECT 0 722.155 0.070 722.785 ;
    RECT 0 722.855 0.070 723.485 ;
    RECT 0 723.555 0.070 724.185 ;
    RECT 0 724.255 0.070 724.885 ;
    RECT 0 724.955 0.070 725.585 ;
    RECT 0 725.655 0.070 726.285 ;
    RECT 0 726.355 0.070 726.985 ;
    RECT 0 727.055 0.070 727.685 ;
    RECT 0 727.755 0.070 728.385 ;
    RECT 0 728.455 0.070 729.085 ;
    RECT 0 729.155 0.070 729.785 ;
    RECT 0 729.855 0.070 730.485 ;
    RECT 0 730.555 0.070 731.185 ;
    RECT 0 731.255 0.070 731.885 ;
    RECT 0 731.955 0.070 732.585 ;
    RECT 0 732.655 0.070 733.285 ;
    RECT 0 733.355 0.070 733.985 ;
    RECT 0 734.055 0.070 734.685 ;
    RECT 0 734.755 0.070 735.385 ;
    RECT 0 735.455 0.070 736.085 ;
    RECT 0 736.155 0.070 736.785 ;
    RECT 0 736.855 0.070 737.485 ;
    RECT 0 737.555 0.070 738.185 ;
    RECT 0 738.255 0.070 738.885 ;
    RECT 0 738.955 0.070 739.585 ;
    RECT 0 739.655 0.070 740.285 ;
    RECT 0 740.355 0.070 740.985 ;
    RECT 0 741.055 0.070 741.685 ;
    RECT 0 741.755 0.070 742.385 ;
    RECT 0 742.455 0.070 743.085 ;
    RECT 0 743.155 0.070 743.785 ;
    RECT 0 743.855 0.070 744.485 ;
    RECT 0 744.555 0.070 745.185 ;
    RECT 0 745.255 0.070 745.885 ;
    RECT 0 745.955 0.070 746.585 ;
    RECT 0 746.655 0.070 747.285 ;
    RECT 0 747.355 0.070 747.985 ;
    RECT 0 748.055 0.070 748.685 ;
    RECT 0 748.755 0.070 749.385 ;
    RECT 0 749.455 0.070 750.085 ;
    RECT 0 750.155 0.070 750.785 ;
    RECT 0 750.855 0.070 751.485 ;
    RECT 0 751.555 0.070 752.185 ;
    RECT 0 752.255 0.070 752.885 ;
    RECT 0 752.955 0.070 753.585 ;
    RECT 0 753.655 0.070 754.285 ;
    RECT 0 754.355 0.070 754.985 ;
    RECT 0 755.055 0.070 755.685 ;
    RECT 0 755.755 0.070 756.385 ;
    RECT 0 756.455 0.070 757.085 ;
    RECT 0 757.155 0.070 757.785 ;
    RECT 0 757.855 0.070 758.485 ;
    RECT 0 758.555 0.070 759.185 ;
    RECT 0 759.255 0.070 759.885 ;
    RECT 0 759.955 0.070 760.585 ;
    RECT 0 760.655 0.070 761.285 ;
    RECT 0 761.355 0.070 761.985 ;
    RECT 0 762.055 0.070 762.685 ;
    RECT 0 762.755 0.070 763.385 ;
    RECT 0 763.455 0.070 764.085 ;
    RECT 0 764.155 0.070 764.785 ;
    RECT 0 764.855 0.070 812.805 ;
    RECT 0 812.875 0.070 813.505 ;
    RECT 0 813.575 0.070 814.205 ;
    RECT 0 814.275 0.070 814.905 ;
    RECT 0 814.975 0.070 815.605 ;
    RECT 0 815.675 0.070 816.305 ;
    RECT 0 816.375 0.070 817.005 ;
    RECT 0 817.075 0.070 817.705 ;
    RECT 0 817.775 0.070 818.405 ;
    RECT 0 818.475 0.070 819.105 ;
    RECT 0 819.175 0.070 819.805 ;
    RECT 0 819.875 0.070 820.505 ;
    RECT 0 820.575 0.070 821.205 ;
    RECT 0 821.275 0.070 821.905 ;
    RECT 0 821.975 0.070 822.605 ;
    RECT 0 822.675 0.070 823.305 ;
    RECT 0 823.375 0.070 824.005 ;
    RECT 0 824.075 0.070 824.705 ;
    RECT 0 824.775 0.070 825.405 ;
    RECT 0 825.475 0.070 826.105 ;
    RECT 0 826.175 0.070 826.805 ;
    RECT 0 826.875 0.070 827.505 ;
    RECT 0 827.575 0.070 828.205 ;
    RECT 0 828.275 0.070 828.905 ;
    RECT 0 828.975 0.070 829.605 ;
    RECT 0 829.675 0.070 830.305 ;
    RECT 0 830.375 0.070 831.005 ;
    RECT 0 831.075 0.070 831.705 ;
    RECT 0 831.775 0.070 832.405 ;
    RECT 0 832.475 0.070 833.105 ;
    RECT 0 833.175 0.070 833.805 ;
    RECT 0 833.875 0.070 834.505 ;
    RECT 0 834.575 0.070 835.205 ;
    RECT 0 835.275 0.070 835.905 ;
    RECT 0 835.975 0.070 836.605 ;
    RECT 0 836.675 0.070 837.305 ;
    RECT 0 837.375 0.070 838.005 ;
    RECT 0 838.075 0.070 838.705 ;
    RECT 0 838.775 0.070 839.405 ;
    RECT 0 839.475 0.070 840.105 ;
    RECT 0 840.175 0.070 840.805 ;
    RECT 0 840.875 0.070 841.505 ;
    RECT 0 841.575 0.070 842.205 ;
    RECT 0 842.275 0.070 842.905 ;
    RECT 0 842.975 0.070 843.605 ;
    RECT 0 843.675 0.070 844.305 ;
    RECT 0 844.375 0.070 845.005 ;
    RECT 0 845.075 0.070 845.705 ;
    RECT 0 845.775 0.070 846.405 ;
    RECT 0 846.475 0.070 847.105 ;
    RECT 0 847.175 0.070 847.805 ;
    RECT 0 847.875 0.070 848.505 ;
    RECT 0 848.575 0.070 849.205 ;
    RECT 0 849.275 0.070 849.905 ;
    RECT 0 849.975 0.070 850.605 ;
    RECT 0 850.675 0.070 851.305 ;
    RECT 0 851.375 0.070 852.005 ;
    RECT 0 852.075 0.070 852.705 ;
    RECT 0 852.775 0.070 853.405 ;
    RECT 0 853.475 0.070 854.105 ;
    RECT 0 854.175 0.070 854.805 ;
    RECT 0 854.875 0.070 855.505 ;
    RECT 0 855.575 0.070 856.205 ;
    RECT 0 856.275 0.070 856.905 ;
    RECT 0 856.975 0.070 857.605 ;
    RECT 0 857.675 0.070 858.305 ;
    RECT 0 858.375 0.070 859.005 ;
    RECT 0 859.075 0.070 859.705 ;
    RECT 0 859.775 0.070 860.405 ;
    RECT 0 860.475 0.070 861.105 ;
    RECT 0 861.175 0.070 861.805 ;
    RECT 0 861.875 0.070 862.505 ;
    RECT 0 862.575 0.070 863.205 ;
    RECT 0 863.275 0.070 863.905 ;
    RECT 0 863.975 0.070 864.605 ;
    RECT 0 864.675 0.070 865.305 ;
    RECT 0 865.375 0.070 866.005 ;
    RECT 0 866.075 0.070 866.705 ;
    RECT 0 866.775 0.070 867.405 ;
    RECT 0 867.475 0.070 868.105 ;
    RECT 0 868.175 0.070 868.805 ;
    RECT 0 868.875 0.070 869.505 ;
    RECT 0 869.575 0.070 870.205 ;
    RECT 0 870.275 0.070 870.905 ;
    RECT 0 870.975 0.070 871.605 ;
    RECT 0 871.675 0.070 872.305 ;
    RECT 0 872.375 0.070 873.005 ;
    RECT 0 873.075 0.070 873.705 ;
    RECT 0 873.775 0.070 874.405 ;
    RECT 0 874.475 0.070 875.105 ;
    RECT 0 875.175 0.070 875.805 ;
    RECT 0 875.875 0.070 876.505 ;
    RECT 0 876.575 0.070 877.205 ;
    RECT 0 877.275 0.070 877.905 ;
    RECT 0 877.975 0.070 878.605 ;
    RECT 0 878.675 0.070 879.305 ;
    RECT 0 879.375 0.070 880.005 ;
    RECT 0 880.075 0.070 880.705 ;
    RECT 0 880.775 0.070 881.405 ;
    RECT 0 881.475 0.070 882.105 ;
    RECT 0 882.175 0.070 882.805 ;
    RECT 0 882.875 0.070 883.505 ;
    RECT 0 883.575 0.070 884.205 ;
    RECT 0 884.275 0.070 884.905 ;
    RECT 0 884.975 0.070 885.605 ;
    RECT 0 885.675 0.070 886.305 ;
    RECT 0 886.375 0.070 887.005 ;
    RECT 0 887.075 0.070 887.705 ;
    RECT 0 887.775 0.070 888.405 ;
    RECT 0 888.475 0.070 889.105 ;
    RECT 0 889.175 0.070 889.805 ;
    RECT 0 889.875 0.070 890.505 ;
    RECT 0 890.575 0.070 891.205 ;
    RECT 0 891.275 0.070 891.905 ;
    RECT 0 891.975 0.070 892.605 ;
    RECT 0 892.675 0.070 893.305 ;
    RECT 0 893.375 0.070 894.005 ;
    RECT 0 894.075 0.070 894.705 ;
    RECT 0 894.775 0.070 895.405 ;
    RECT 0 895.475 0.070 896.105 ;
    RECT 0 896.175 0.070 896.805 ;
    RECT 0 896.875 0.070 897.505 ;
    RECT 0 897.575 0.070 898.205 ;
    RECT 0 898.275 0.070 898.905 ;
    RECT 0 898.975 0.070 899.605 ;
    RECT 0 899.675 0.070 900.305 ;
    RECT 0 900.375 0.070 901.005 ;
    RECT 0 901.075 0.070 901.705 ;
    RECT 0 901.775 0.070 902.405 ;
    RECT 0 902.475 0.070 903.105 ;
    RECT 0 903.175 0.070 903.805 ;
    RECT 0 903.875 0.070 904.505 ;
    RECT 0 904.575 0.070 905.205 ;
    RECT 0 905.275 0.070 905.905 ;
    RECT 0 905.975 0.070 906.605 ;
    RECT 0 906.675 0.070 907.305 ;
    RECT 0 907.375 0.070 908.005 ;
    RECT 0 908.075 0.070 908.705 ;
    RECT 0 908.775 0.070 909.405 ;
    RECT 0 909.475 0.070 910.105 ;
    RECT 0 910.175 0.070 910.805 ;
    RECT 0 910.875 0.070 911.505 ;
    RECT 0 911.575 0.070 912.205 ;
    RECT 0 912.275 0.070 912.905 ;
    RECT 0 912.975 0.070 913.605 ;
    RECT 0 913.675 0.070 914.305 ;
    RECT 0 914.375 0.070 915.005 ;
    RECT 0 915.075 0.070 915.705 ;
    RECT 0 915.775 0.070 916.405 ;
    RECT 0 916.475 0.070 917.105 ;
    RECT 0 917.175 0.070 917.805 ;
    RECT 0 917.875 0.070 918.505 ;
    RECT 0 918.575 0.070 919.205 ;
    RECT 0 919.275 0.070 919.905 ;
    RECT 0 919.975 0.070 920.605 ;
    RECT 0 920.675 0.070 921.305 ;
    RECT 0 921.375 0.070 922.005 ;
    RECT 0 922.075 0.070 922.705 ;
    RECT 0 922.775 0.070 923.405 ;
    RECT 0 923.475 0.070 924.105 ;
    RECT 0 924.175 0.070 924.805 ;
    RECT 0 924.875 0.070 925.505 ;
    RECT 0 925.575 0.070 926.205 ;
    RECT 0 926.275 0.070 926.905 ;
    RECT 0 926.975 0.070 927.605 ;
    RECT 0 927.675 0.070 928.305 ;
    RECT 0 928.375 0.070 929.005 ;
    RECT 0 929.075 0.070 929.705 ;
    RECT 0 929.775 0.070 930.405 ;
    RECT 0 930.475 0.070 931.105 ;
    RECT 0 931.175 0.070 931.805 ;
    RECT 0 931.875 0.070 932.505 ;
    RECT 0 932.575 0.070 933.205 ;
    RECT 0 933.275 0.070 933.905 ;
    RECT 0 933.975 0.070 934.605 ;
    RECT 0 934.675 0.070 935.305 ;
    RECT 0 935.375 0.070 936.005 ;
    RECT 0 936.075 0.070 936.705 ;
    RECT 0 936.775 0.070 937.405 ;
    RECT 0 937.475 0.070 938.105 ;
    RECT 0 938.175 0.070 938.805 ;
    RECT 0 938.875 0.070 939.505 ;
    RECT 0 939.575 0.070 940.205 ;
    RECT 0 940.275 0.070 940.905 ;
    RECT 0 940.975 0.070 941.605 ;
    RECT 0 941.675 0.070 942.305 ;
    RECT 0 942.375 0.070 943.005 ;
    RECT 0 943.075 0.070 943.705 ;
    RECT 0 943.775 0.070 944.405 ;
    RECT 0 944.475 0.070 945.105 ;
    RECT 0 945.175 0.070 945.805 ;
    RECT 0 945.875 0.070 946.505 ;
    RECT 0 946.575 0.070 947.205 ;
    RECT 0 947.275 0.070 947.905 ;
    RECT 0 947.975 0.070 948.605 ;
    RECT 0 948.675 0.070 949.305 ;
    RECT 0 949.375 0.070 950.005 ;
    RECT 0 950.075 0.070 950.705 ;
    RECT 0 950.775 0.070 951.405 ;
    RECT 0 951.475 0.070 952.105 ;
    RECT 0 952.175 0.070 952.805 ;
    RECT 0 952.875 0.070 953.505 ;
    RECT 0 953.575 0.070 954.205 ;
    RECT 0 954.275 0.070 954.905 ;
    RECT 0 954.975 0.070 955.605 ;
    RECT 0 955.675 0.070 956.305 ;
    RECT 0 956.375 0.070 957.005 ;
    RECT 0 957.075 0.070 957.705 ;
    RECT 0 957.775 0.070 958.405 ;
    RECT 0 958.475 0.070 959.105 ;
    RECT 0 959.175 0.070 959.805 ;
    RECT 0 959.875 0.070 960.505 ;
    RECT 0 960.575 0.070 961.205 ;
    RECT 0 961.275 0.070 961.905 ;
    RECT 0 961.975 0.070 962.605 ;
    RECT 0 962.675 0.070 963.305 ;
    RECT 0 963.375 0.070 964.005 ;
    RECT 0 964.075 0.070 964.705 ;
    RECT 0 964.775 0.070 965.405 ;
    RECT 0 965.475 0.070 966.105 ;
    RECT 0 966.175 0.070 966.805 ;
    RECT 0 966.875 0.070 967.505 ;
    RECT 0 967.575 0.070 968.205 ;
    RECT 0 968.275 0.070 968.905 ;
    RECT 0 968.975 0.070 969.605 ;
    RECT 0 969.675 0.070 970.305 ;
    RECT 0 970.375 0.070 971.005 ;
    RECT 0 971.075 0.070 971.705 ;
    RECT 0 971.775 0.070 972.405 ;
    RECT 0 972.475 0.070 973.105 ;
    RECT 0 973.175 0.070 973.805 ;
    RECT 0 973.875 0.070 974.505 ;
    RECT 0 974.575 0.070 975.205 ;
    RECT 0 975.275 0.070 975.905 ;
    RECT 0 975.975 0.070 976.605 ;
    RECT 0 976.675 0.070 977.305 ;
    RECT 0 977.375 0.070 978.005 ;
    RECT 0 978.075 0.070 978.705 ;
    RECT 0 978.775 0.070 979.405 ;
    RECT 0 979.475 0.070 980.105 ;
    RECT 0 980.175 0.070 980.805 ;
    RECT 0 980.875 0.070 981.505 ;
    RECT 0 981.575 0.070 982.205 ;
    RECT 0 982.275 0.070 982.905 ;
    RECT 0 982.975 0.070 983.605 ;
    RECT 0 983.675 0.070 984.305 ;
    RECT 0 984.375 0.070 985.005 ;
    RECT 0 985.075 0.070 985.705 ;
    RECT 0 985.775 0.070 986.405 ;
    RECT 0 986.475 0.070 987.105 ;
    RECT 0 987.175 0.070 987.805 ;
    RECT 0 987.875 0.070 988.505 ;
    RECT 0 988.575 0.070 989.205 ;
    RECT 0 989.275 0.070 989.905 ;
    RECT 0 989.975 0.070 990.605 ;
    RECT 0 990.675 0.070 991.305 ;
    RECT 0 991.375 0.070 992.005 ;
    RECT 0 992.075 0.070 992.705 ;
    RECT 0 992.775 0.070 993.405 ;
    RECT 0 993.475 0.070 994.105 ;
    RECT 0 994.175 0.070 994.805 ;
    RECT 0 994.875 0.070 995.505 ;
    RECT 0 995.575 0.070 996.205 ;
    RECT 0 996.275 0.070 996.905 ;
    RECT 0 996.975 0.070 997.605 ;
    RECT 0 997.675 0.070 998.305 ;
    RECT 0 998.375 0.070 999.005 ;
    RECT 0 999.075 0.070 999.705 ;
    RECT 0 999.775 0.070 1000.405 ;
    RECT 0 1000.475 0.070 1001.105 ;
    RECT 0 1001.175 0.070 1001.805 ;
    RECT 0 1001.875 0.070 1002.505 ;
    RECT 0 1002.575 0.070 1003.205 ;
    RECT 0 1003.275 0.070 1003.905 ;
    RECT 0 1003.975 0.070 1004.605 ;
    RECT 0 1004.675 0.070 1005.305 ;
    RECT 0 1005.375 0.070 1006.005 ;
    RECT 0 1006.075 0.070 1006.705 ;
    RECT 0 1006.775 0.070 1007.405 ;
    RECT 0 1007.475 0.070 1008.105 ;
    RECT 0 1008.175 0.070 1008.805 ;
    RECT 0 1008.875 0.070 1009.505 ;
    RECT 0 1009.575 0.070 1010.205 ;
    RECT 0 1010.275 0.070 1010.905 ;
    RECT 0 1010.975 0.070 1011.605 ;
    RECT 0 1011.675 0.070 1012.305 ;
    RECT 0 1012.375 0.070 1013.005 ;
    RECT 0 1013.075 0.070 1013.705 ;
    RECT 0 1013.775 0.070 1014.405 ;
    RECT 0 1014.475 0.070 1015.105 ;
    RECT 0 1015.175 0.070 1015.805 ;
    RECT 0 1015.875 0.070 1016.505 ;
    RECT 0 1016.575 0.070 1017.205 ;
    RECT 0 1017.275 0.070 1017.905 ;
    RECT 0 1017.975 0.070 1018.605 ;
    RECT 0 1018.675 0.070 1019.305 ;
    RECT 0 1019.375 0.070 1020.005 ;
    RECT 0 1020.075 0.070 1020.705 ;
    RECT 0 1020.775 0.070 1021.405 ;
    RECT 0 1021.475 0.070 1022.105 ;
    RECT 0 1022.175 0.070 1022.805 ;
    RECT 0 1022.875 0.070 1023.505 ;
    RECT 0 1023.575 0.070 1024.205 ;
    RECT 0 1024.275 0.070 1024.905 ;
    RECT 0 1024.975 0.070 1025.605 ;
    RECT 0 1025.675 0.070 1026.305 ;
    RECT 0 1026.375 0.070 1027.005 ;
    RECT 0 1027.075 0.070 1027.705 ;
    RECT 0 1027.775 0.070 1028.405 ;
    RECT 0 1028.475 0.070 1029.105 ;
    RECT 0 1029.175 0.070 1029.805 ;
    RECT 0 1029.875 0.070 1030.505 ;
    RECT 0 1030.575 0.070 1031.205 ;
    RECT 0 1031.275 0.070 1031.905 ;
    RECT 0 1031.975 0.070 1032.605 ;
    RECT 0 1032.675 0.070 1033.305 ;
    RECT 0 1033.375 0.070 1034.005 ;
    RECT 0 1034.075 0.070 1034.705 ;
    RECT 0 1034.775 0.070 1035.405 ;
    RECT 0 1035.475 0.070 1036.105 ;
    RECT 0 1036.175 0.070 1036.805 ;
    RECT 0 1036.875 0.070 1037.505 ;
    RECT 0 1037.575 0.070 1038.205 ;
    RECT 0 1038.275 0.070 1038.905 ;
    RECT 0 1038.975 0.070 1039.605 ;
    RECT 0 1039.675 0.070 1040.305 ;
    RECT 0 1040.375 0.070 1041.005 ;
    RECT 0 1041.075 0.070 1041.705 ;
    RECT 0 1041.775 0.070 1042.405 ;
    RECT 0 1042.475 0.070 1043.105 ;
    RECT 0 1043.175 0.070 1043.805 ;
    RECT 0 1043.875 0.070 1044.505 ;
    RECT 0 1044.575 0.070 1045.205 ;
    RECT 0 1045.275 0.070 1045.905 ;
    RECT 0 1045.975 0.070 1046.605 ;
    RECT 0 1046.675 0.070 1047.305 ;
    RECT 0 1047.375 0.070 1048.005 ;
    RECT 0 1048.075 0.070 1048.705 ;
    RECT 0 1048.775 0.070 1049.405 ;
    RECT 0 1049.475 0.070 1050.105 ;
    RECT 0 1050.175 0.070 1050.805 ;
    RECT 0 1050.875 0.070 1051.505 ;
    RECT 0 1051.575 0.070 1052.205 ;
    RECT 0 1052.275 0.070 1052.905 ;
    RECT 0 1052.975 0.070 1053.605 ;
    RECT 0 1053.675 0.070 1054.305 ;
    RECT 0 1054.375 0.070 1055.005 ;
    RECT 0 1055.075 0.070 1055.705 ;
    RECT 0 1055.775 0.070 1056.405 ;
    RECT 0 1056.475 0.070 1057.105 ;
    RECT 0 1057.175 0.070 1057.805 ;
    RECT 0 1057.875 0.070 1058.505 ;
    RECT 0 1058.575 0.070 1059.205 ;
    RECT 0 1059.275 0.070 1059.905 ;
    RECT 0 1059.975 0.070 1060.605 ;
    RECT 0 1060.675 0.070 1061.305 ;
    RECT 0 1061.375 0.070 1062.005 ;
    RECT 0 1062.075 0.070 1062.705 ;
    RECT 0 1062.775 0.070 1063.405 ;
    RECT 0 1063.475 0.070 1064.105 ;
    RECT 0 1064.175 0.070 1064.805 ;
    RECT 0 1064.875 0.070 1065.505 ;
    RECT 0 1065.575 0.070 1066.205 ;
    RECT 0 1066.275 0.070 1066.905 ;
    RECT 0 1066.975 0.070 1067.605 ;
    RECT 0 1067.675 0.070 1068.305 ;
    RECT 0 1068.375 0.070 1069.005 ;
    RECT 0 1069.075 0.070 1069.705 ;
    RECT 0 1069.775 0.070 1070.405 ;
    RECT 0 1070.475 0.070 1071.105 ;
    RECT 0 1071.175 0.070 1071.805 ;
    RECT 0 1071.875 0.070 1072.505 ;
    RECT 0 1072.575 0.070 1073.205 ;
    RECT 0 1073.275 0.070 1073.905 ;
    RECT 0 1073.975 0.070 1074.605 ;
    RECT 0 1074.675 0.070 1075.305 ;
    RECT 0 1075.375 0.070 1076.005 ;
    RECT 0 1076.075 0.070 1076.705 ;
    RECT 0 1076.775 0.070 1077.405 ;
    RECT 0 1077.475 0.070 1078.105 ;
    RECT 0 1078.175 0.070 1078.805 ;
    RECT 0 1078.875 0.070 1079.505 ;
    RECT 0 1079.575 0.070 1080.205 ;
    RECT 0 1080.275 0.070 1080.905 ;
    RECT 0 1080.975 0.070 1081.605 ;
    RECT 0 1081.675 0.070 1082.305 ;
    RECT 0 1082.375 0.070 1083.005 ;
    RECT 0 1083.075 0.070 1083.705 ;
    RECT 0 1083.775 0.070 1084.405 ;
    RECT 0 1084.475 0.070 1085.105 ;
    RECT 0 1085.175 0.070 1085.805 ;
    RECT 0 1085.875 0.070 1086.505 ;
    RECT 0 1086.575 0.070 1087.205 ;
    RECT 0 1087.275 0.070 1087.905 ;
    RECT 0 1087.975 0.070 1088.605 ;
    RECT 0 1088.675 0.070 1089.305 ;
    RECT 0 1089.375 0.070 1090.005 ;
    RECT 0 1090.075 0.070 1090.705 ;
    RECT 0 1090.775 0.070 1091.405 ;
    RECT 0 1091.475 0.070 1092.105 ;
    RECT 0 1092.175 0.070 1092.805 ;
    RECT 0 1092.875 0.070 1093.505 ;
    RECT 0 1093.575 0.070 1094.205 ;
    RECT 0 1094.275 0.070 1094.905 ;
    RECT 0 1094.975 0.070 1095.605 ;
    RECT 0 1095.675 0.070 1096.305 ;
    RECT 0 1096.375 0.070 1097.005 ;
    RECT 0 1097.075 0.070 1097.705 ;
    RECT 0 1097.775 0.070 1098.405 ;
    RECT 0 1098.475 0.070 1099.105 ;
    RECT 0 1099.175 0.070 1099.805 ;
    RECT 0 1099.875 0.070 1100.505 ;
    RECT 0 1100.575 0.070 1101.205 ;
    RECT 0 1101.275 0.070 1101.905 ;
    RECT 0 1101.975 0.070 1102.605 ;
    RECT 0 1102.675 0.070 1103.305 ;
    RECT 0 1103.375 0.070 1104.005 ;
    RECT 0 1104.075 0.070 1104.705 ;
    RECT 0 1104.775 0.070 1105.405 ;
    RECT 0 1105.475 0.070 1106.105 ;
    RECT 0 1106.175 0.070 1106.805 ;
    RECT 0 1106.875 0.070 1107.505 ;
    RECT 0 1107.575 0.070 1108.205 ;
    RECT 0 1108.275 0.070 1108.905 ;
    RECT 0 1108.975 0.070 1109.605 ;
    RECT 0 1109.675 0.070 1110.305 ;
    RECT 0 1110.375 0.070 1111.005 ;
    RECT 0 1111.075 0.070 1111.705 ;
    RECT 0 1111.775 0.070 1112.405 ;
    RECT 0 1112.475 0.070 1113.105 ;
    RECT 0 1113.175 0.070 1113.805 ;
    RECT 0 1113.875 0.070 1114.505 ;
    RECT 0 1114.575 0.070 1115.205 ;
    RECT 0 1115.275 0.070 1115.905 ;
    RECT 0 1115.975 0.070 1116.605 ;
    RECT 0 1116.675 0.070 1117.305 ;
    RECT 0 1117.375 0.070 1118.005 ;
    RECT 0 1118.075 0.070 1118.705 ;
    RECT 0 1118.775 0.070 1119.405 ;
    RECT 0 1119.475 0.070 1120.105 ;
    RECT 0 1120.175 0.070 1120.805 ;
    RECT 0 1120.875 0.070 1121.505 ;
    RECT 0 1121.575 0.070 1122.205 ;
    RECT 0 1122.275 0.070 1122.905 ;
    RECT 0 1122.975 0.070 1123.605 ;
    RECT 0 1123.675 0.070 1124.305 ;
    RECT 0 1124.375 0.070 1125.005 ;
    RECT 0 1125.075 0.070 1125.705 ;
    RECT 0 1125.775 0.070 1126.405 ;
    RECT 0 1126.475 0.070 1127.105 ;
    RECT 0 1127.175 0.070 1127.805 ;
    RECT 0 1127.875 0.070 1128.505 ;
    RECT 0 1128.575 0.070 1129.205 ;
    RECT 0 1129.275 0.070 1129.905 ;
    RECT 0 1129.975 0.070 1130.605 ;
    RECT 0 1130.675 0.070 1131.305 ;
    RECT 0 1131.375 0.070 1132.005 ;
    RECT 0 1132.075 0.070 1132.705 ;
    RECT 0 1132.775 0.070 1133.405 ;
    RECT 0 1133.475 0.070 1134.105 ;
    RECT 0 1134.175 0.070 1134.805 ;
    RECT 0 1134.875 0.070 1135.505 ;
    RECT 0 1135.575 0.070 1136.205 ;
    RECT 0 1136.275 0.070 1136.905 ;
    RECT 0 1136.975 0.070 1137.605 ;
    RECT 0 1137.675 0.070 1138.305 ;
    RECT 0 1138.375 0.070 1139.005 ;
    RECT 0 1139.075 0.070 1139.705 ;
    RECT 0 1139.775 0.070 1140.405 ;
    RECT 0 1140.475 0.070 1141.105 ;
    RECT 0 1141.175 0.070 1141.805 ;
    RECT 0 1141.875 0.070 1142.505 ;
    RECT 0 1142.575 0.070 1143.205 ;
    RECT 0 1143.275 0.070 1143.905 ;
    RECT 0 1143.975 0.070 1144.605 ;
    RECT 0 1144.675 0.070 1145.305 ;
    RECT 0 1145.375 0.070 1146.005 ;
    RECT 0 1146.075 0.070 1146.705 ;
    RECT 0 1146.775 0.070 1147.405 ;
    RECT 0 1147.475 0.070 1148.105 ;
    RECT 0 1148.175 0.070 1148.805 ;
    RECT 0 1148.875 0.070 1149.505 ;
    RECT 0 1149.575 0.070 1150.205 ;
    RECT 0 1150.275 0.070 1150.905 ;
    RECT 0 1150.975 0.070 1151.605 ;
    RECT 0 1151.675 0.070 1152.305 ;
    RECT 0 1152.375 0.070 1153.005 ;
    RECT 0 1153.075 0.070 1153.705 ;
    RECT 0 1153.775 0.070 1154.405 ;
    RECT 0 1154.475 0.070 1155.105 ;
    RECT 0 1155.175 0.070 1155.805 ;
    RECT 0 1155.875 0.070 1156.505 ;
    RECT 0 1156.575 0.070 1157.205 ;
    RECT 0 1157.275 0.070 1157.905 ;
    RECT 0 1157.975 0.070 1158.605 ;
    RECT 0 1158.675 0.070 1159.305 ;
    RECT 0 1159.375 0.070 1160.005 ;
    RECT 0 1160.075 0.070 1160.705 ;
    RECT 0 1160.775 0.070 1161.405 ;
    RECT 0 1161.475 0.070 1162.105 ;
    RECT 0 1162.175 0.070 1162.805 ;
    RECT 0 1162.875 0.070 1163.505 ;
    RECT 0 1163.575 0.070 1164.205 ;
    RECT 0 1164.275 0.070 1164.905 ;
    RECT 0 1164.975 0.070 1165.605 ;
    RECT 0 1165.675 0.070 1166.305 ;
    RECT 0 1166.375 0.070 1167.005 ;
    RECT 0 1167.075 0.070 1167.705 ;
    RECT 0 1167.775 0.070 1168.405 ;
    RECT 0 1168.475 0.070 1169.105 ;
    RECT 0 1169.175 0.070 1169.805 ;
    RECT 0 1169.875 0.070 1170.505 ;
    RECT 0 1170.575 0.070 1218.525 ;
    RECT 0 1218.595 0.070 1219.225 ;
    RECT 0 1219.295 0.070 1219.925 ;
    RECT 0 1219.995 0.070 1220.625 ;
    RECT 0 1220.695 0.070 1221.325 ;
    RECT 0 1221.395 0.070 1222.025 ;
    RECT 0 1222.095 0.070 1222.725 ;
    RECT 0 1222.795 0.070 1223.425 ;
    RECT 0 1223.495 0.070 1224.125 ;
    RECT 0 1224.195 0.070 1224.825 ;
    RECT 0 1224.895 0.070 1225.525 ;
    RECT 0 1225.595 0.070 1226.225 ;
    RECT 0 1226.295 0.070 1274.245 ;
    RECT 0 1274.315 0.070 1274.945 ;
    RECT 0 1275.015 0.070 1275.645 ;
    RECT 0 1275.715 0.070 1281.000 ;
    LAYER metal4 ;
    RECT 0 0 2064.540 1.400 ;
    RECT 0 1279.600 2064.540 1281.000 ;
    RECT 0.000 1.400 1.260 1279.600 ;
    RECT 1.540 1.400 2.380 1279.600 ;
    RECT 2.660 1.400 3.500 1279.600 ;
    RECT 3.780 1.400 4.620 1279.600 ;
    RECT 4.900 1.400 5.740 1279.600 ;
    RECT 6.020 1.400 6.860 1279.600 ;
    RECT 7.140 1.400 7.980 1279.600 ;
    RECT 8.260 1.400 9.100 1279.600 ;
    RECT 9.380 1.400 10.220 1279.600 ;
    RECT 10.500 1.400 11.340 1279.600 ;
    RECT 11.620 1.400 12.460 1279.600 ;
    RECT 12.740 1.400 13.580 1279.600 ;
    RECT 13.860 1.400 14.700 1279.600 ;
    RECT 14.980 1.400 15.820 1279.600 ;
    RECT 16.100 1.400 16.940 1279.600 ;
    RECT 17.220 1.400 18.060 1279.600 ;
    RECT 18.340 1.400 19.180 1279.600 ;
    RECT 19.460 1.400 20.300 1279.600 ;
    RECT 20.580 1.400 21.420 1279.600 ;
    RECT 21.700 1.400 22.540 1279.600 ;
    RECT 22.820 1.400 23.660 1279.600 ;
    RECT 23.940 1.400 24.780 1279.600 ;
    RECT 25.060 1.400 25.900 1279.600 ;
    RECT 26.180 1.400 27.020 1279.600 ;
    RECT 27.300 1.400 28.140 1279.600 ;
    RECT 28.420 1.400 29.260 1279.600 ;
    RECT 29.540 1.400 30.380 1279.600 ;
    RECT 30.660 1.400 31.500 1279.600 ;
    RECT 31.780 1.400 32.620 1279.600 ;
    RECT 32.900 1.400 33.740 1279.600 ;
    RECT 34.020 1.400 34.860 1279.600 ;
    RECT 35.140 1.400 35.980 1279.600 ;
    RECT 36.260 1.400 37.100 1279.600 ;
    RECT 37.380 1.400 38.220 1279.600 ;
    RECT 38.500 1.400 39.340 1279.600 ;
    RECT 39.620 1.400 40.460 1279.600 ;
    RECT 40.740 1.400 41.580 1279.600 ;
    RECT 41.860 1.400 42.700 1279.600 ;
    RECT 42.980 1.400 43.820 1279.600 ;
    RECT 44.100 1.400 44.940 1279.600 ;
    RECT 45.220 1.400 46.060 1279.600 ;
    RECT 46.340 1.400 47.180 1279.600 ;
    RECT 47.460 1.400 48.300 1279.600 ;
    RECT 48.580 1.400 49.420 1279.600 ;
    RECT 49.700 1.400 50.540 1279.600 ;
    RECT 50.820 1.400 51.660 1279.600 ;
    RECT 51.940 1.400 52.780 1279.600 ;
    RECT 53.060 1.400 53.900 1279.600 ;
    RECT 54.180 1.400 55.020 1279.600 ;
    RECT 55.300 1.400 56.140 1279.600 ;
    RECT 56.420 1.400 57.260 1279.600 ;
    RECT 57.540 1.400 58.380 1279.600 ;
    RECT 58.660 1.400 59.500 1279.600 ;
    RECT 59.780 1.400 60.620 1279.600 ;
    RECT 60.900 1.400 61.740 1279.600 ;
    RECT 62.020 1.400 62.860 1279.600 ;
    RECT 63.140 1.400 63.980 1279.600 ;
    RECT 64.260 1.400 65.100 1279.600 ;
    RECT 65.380 1.400 66.220 1279.600 ;
    RECT 66.500 1.400 67.340 1279.600 ;
    RECT 67.620 1.400 68.460 1279.600 ;
    RECT 68.740 1.400 69.580 1279.600 ;
    RECT 69.860 1.400 70.700 1279.600 ;
    RECT 70.980 1.400 71.820 1279.600 ;
    RECT 72.100 1.400 72.940 1279.600 ;
    RECT 73.220 1.400 74.060 1279.600 ;
    RECT 74.340 1.400 75.180 1279.600 ;
    RECT 75.460 1.400 76.300 1279.600 ;
    RECT 76.580 1.400 77.420 1279.600 ;
    RECT 77.700 1.400 78.540 1279.600 ;
    RECT 78.820 1.400 79.660 1279.600 ;
    RECT 79.940 1.400 80.780 1279.600 ;
    RECT 81.060 1.400 81.900 1279.600 ;
    RECT 82.180 1.400 83.020 1279.600 ;
    RECT 83.300 1.400 84.140 1279.600 ;
    RECT 84.420 1.400 85.260 1279.600 ;
    RECT 85.540 1.400 86.380 1279.600 ;
    RECT 86.660 1.400 87.500 1279.600 ;
    RECT 87.780 1.400 88.620 1279.600 ;
    RECT 88.900 1.400 89.740 1279.600 ;
    RECT 90.020 1.400 90.860 1279.600 ;
    RECT 91.140 1.400 91.980 1279.600 ;
    RECT 92.260 1.400 93.100 1279.600 ;
    RECT 93.380 1.400 94.220 1279.600 ;
    RECT 94.500 1.400 95.340 1279.600 ;
    RECT 95.620 1.400 96.460 1279.600 ;
    RECT 96.740 1.400 97.580 1279.600 ;
    RECT 97.860 1.400 98.700 1279.600 ;
    RECT 98.980 1.400 99.820 1279.600 ;
    RECT 100.100 1.400 100.940 1279.600 ;
    RECT 101.220 1.400 102.060 1279.600 ;
    RECT 102.340 1.400 103.180 1279.600 ;
    RECT 103.460 1.400 104.300 1279.600 ;
    RECT 104.580 1.400 105.420 1279.600 ;
    RECT 105.700 1.400 106.540 1279.600 ;
    RECT 106.820 1.400 107.660 1279.600 ;
    RECT 107.940 1.400 108.780 1279.600 ;
    RECT 109.060 1.400 109.900 1279.600 ;
    RECT 110.180 1.400 111.020 1279.600 ;
    RECT 111.300 1.400 112.140 1279.600 ;
    RECT 112.420 1.400 113.260 1279.600 ;
    RECT 113.540 1.400 114.380 1279.600 ;
    RECT 114.660 1.400 115.500 1279.600 ;
    RECT 115.780 1.400 116.620 1279.600 ;
    RECT 116.900 1.400 117.740 1279.600 ;
    RECT 118.020 1.400 118.860 1279.600 ;
    RECT 119.140 1.400 119.980 1279.600 ;
    RECT 120.260 1.400 121.100 1279.600 ;
    RECT 121.380 1.400 122.220 1279.600 ;
    RECT 122.500 1.400 123.340 1279.600 ;
    RECT 123.620 1.400 124.460 1279.600 ;
    RECT 124.740 1.400 125.580 1279.600 ;
    RECT 125.860 1.400 126.700 1279.600 ;
    RECT 126.980 1.400 127.820 1279.600 ;
    RECT 128.100 1.400 128.940 1279.600 ;
    RECT 129.220 1.400 130.060 1279.600 ;
    RECT 130.340 1.400 131.180 1279.600 ;
    RECT 131.460 1.400 132.300 1279.600 ;
    RECT 132.580 1.400 133.420 1279.600 ;
    RECT 133.700 1.400 134.540 1279.600 ;
    RECT 134.820 1.400 135.660 1279.600 ;
    RECT 135.940 1.400 136.780 1279.600 ;
    RECT 137.060 1.400 137.900 1279.600 ;
    RECT 138.180 1.400 139.020 1279.600 ;
    RECT 139.300 1.400 140.140 1279.600 ;
    RECT 140.420 1.400 141.260 1279.600 ;
    RECT 141.540 1.400 142.380 1279.600 ;
    RECT 142.660 1.400 143.500 1279.600 ;
    RECT 143.780 1.400 144.620 1279.600 ;
    RECT 144.900 1.400 145.740 1279.600 ;
    RECT 146.020 1.400 146.860 1279.600 ;
    RECT 147.140 1.400 147.980 1279.600 ;
    RECT 148.260 1.400 149.100 1279.600 ;
    RECT 149.380 1.400 150.220 1279.600 ;
    RECT 150.500 1.400 151.340 1279.600 ;
    RECT 151.620 1.400 152.460 1279.600 ;
    RECT 152.740 1.400 153.580 1279.600 ;
    RECT 153.860 1.400 154.700 1279.600 ;
    RECT 154.980 1.400 155.820 1279.600 ;
    RECT 156.100 1.400 156.940 1279.600 ;
    RECT 157.220 1.400 158.060 1279.600 ;
    RECT 158.340 1.400 159.180 1279.600 ;
    RECT 159.460 1.400 160.300 1279.600 ;
    RECT 160.580 1.400 161.420 1279.600 ;
    RECT 161.700 1.400 162.540 1279.600 ;
    RECT 162.820 1.400 163.660 1279.600 ;
    RECT 163.940 1.400 164.780 1279.600 ;
    RECT 165.060 1.400 165.900 1279.600 ;
    RECT 166.180 1.400 167.020 1279.600 ;
    RECT 167.300 1.400 168.140 1279.600 ;
    RECT 168.420 1.400 169.260 1279.600 ;
    RECT 169.540 1.400 170.380 1279.600 ;
    RECT 170.660 1.400 171.500 1279.600 ;
    RECT 171.780 1.400 172.620 1279.600 ;
    RECT 172.900 1.400 173.740 1279.600 ;
    RECT 174.020 1.400 174.860 1279.600 ;
    RECT 175.140 1.400 175.980 1279.600 ;
    RECT 176.260 1.400 177.100 1279.600 ;
    RECT 177.380 1.400 178.220 1279.600 ;
    RECT 178.500 1.400 179.340 1279.600 ;
    RECT 179.620 1.400 180.460 1279.600 ;
    RECT 180.740 1.400 181.580 1279.600 ;
    RECT 181.860 1.400 182.700 1279.600 ;
    RECT 182.980 1.400 183.820 1279.600 ;
    RECT 184.100 1.400 184.940 1279.600 ;
    RECT 185.220 1.400 186.060 1279.600 ;
    RECT 186.340 1.400 187.180 1279.600 ;
    RECT 187.460 1.400 188.300 1279.600 ;
    RECT 188.580 1.400 189.420 1279.600 ;
    RECT 189.700 1.400 190.540 1279.600 ;
    RECT 190.820 1.400 191.660 1279.600 ;
    RECT 191.940 1.400 192.780 1279.600 ;
    RECT 193.060 1.400 193.900 1279.600 ;
    RECT 194.180 1.400 195.020 1279.600 ;
    RECT 195.300 1.400 196.140 1279.600 ;
    RECT 196.420 1.400 197.260 1279.600 ;
    RECT 197.540 1.400 198.380 1279.600 ;
    RECT 198.660 1.400 199.500 1279.600 ;
    RECT 199.780 1.400 200.620 1279.600 ;
    RECT 200.900 1.400 201.740 1279.600 ;
    RECT 202.020 1.400 202.860 1279.600 ;
    RECT 203.140 1.400 203.980 1279.600 ;
    RECT 204.260 1.400 205.100 1279.600 ;
    RECT 205.380 1.400 206.220 1279.600 ;
    RECT 206.500 1.400 207.340 1279.600 ;
    RECT 207.620 1.400 208.460 1279.600 ;
    RECT 208.740 1.400 209.580 1279.600 ;
    RECT 209.860 1.400 210.700 1279.600 ;
    RECT 210.980 1.400 211.820 1279.600 ;
    RECT 212.100 1.400 212.940 1279.600 ;
    RECT 213.220 1.400 214.060 1279.600 ;
    RECT 214.340 1.400 215.180 1279.600 ;
    RECT 215.460 1.400 216.300 1279.600 ;
    RECT 216.580 1.400 217.420 1279.600 ;
    RECT 217.700 1.400 218.540 1279.600 ;
    RECT 218.820 1.400 219.660 1279.600 ;
    RECT 219.940 1.400 220.780 1279.600 ;
    RECT 221.060 1.400 221.900 1279.600 ;
    RECT 222.180 1.400 223.020 1279.600 ;
    RECT 223.300 1.400 224.140 1279.600 ;
    RECT 224.420 1.400 225.260 1279.600 ;
    RECT 225.540 1.400 226.380 1279.600 ;
    RECT 226.660 1.400 227.500 1279.600 ;
    RECT 227.780 1.400 228.620 1279.600 ;
    RECT 228.900 1.400 229.740 1279.600 ;
    RECT 230.020 1.400 230.860 1279.600 ;
    RECT 231.140 1.400 231.980 1279.600 ;
    RECT 232.260 1.400 233.100 1279.600 ;
    RECT 233.380 1.400 234.220 1279.600 ;
    RECT 234.500 1.400 235.340 1279.600 ;
    RECT 235.620 1.400 236.460 1279.600 ;
    RECT 236.740 1.400 237.580 1279.600 ;
    RECT 237.860 1.400 238.700 1279.600 ;
    RECT 238.980 1.400 239.820 1279.600 ;
    RECT 240.100 1.400 240.940 1279.600 ;
    RECT 241.220 1.400 242.060 1279.600 ;
    RECT 242.340 1.400 243.180 1279.600 ;
    RECT 243.460 1.400 244.300 1279.600 ;
    RECT 244.580 1.400 245.420 1279.600 ;
    RECT 245.700 1.400 246.540 1279.600 ;
    RECT 246.820 1.400 247.660 1279.600 ;
    RECT 247.940 1.400 248.780 1279.600 ;
    RECT 249.060 1.400 249.900 1279.600 ;
    RECT 250.180 1.400 251.020 1279.600 ;
    RECT 251.300 1.400 252.140 1279.600 ;
    RECT 252.420 1.400 253.260 1279.600 ;
    RECT 253.540 1.400 254.380 1279.600 ;
    RECT 254.660 1.400 255.500 1279.600 ;
    RECT 255.780 1.400 256.620 1279.600 ;
    RECT 256.900 1.400 257.740 1279.600 ;
    RECT 258.020 1.400 258.860 1279.600 ;
    RECT 259.140 1.400 259.980 1279.600 ;
    RECT 260.260 1.400 261.100 1279.600 ;
    RECT 261.380 1.400 262.220 1279.600 ;
    RECT 262.500 1.400 263.340 1279.600 ;
    RECT 263.620 1.400 264.460 1279.600 ;
    RECT 264.740 1.400 265.580 1279.600 ;
    RECT 265.860 1.400 266.700 1279.600 ;
    RECT 266.980 1.400 267.820 1279.600 ;
    RECT 268.100 1.400 268.940 1279.600 ;
    RECT 269.220 1.400 270.060 1279.600 ;
    RECT 270.340 1.400 271.180 1279.600 ;
    RECT 271.460 1.400 272.300 1279.600 ;
    RECT 272.580 1.400 273.420 1279.600 ;
    RECT 273.700 1.400 274.540 1279.600 ;
    RECT 274.820 1.400 275.660 1279.600 ;
    RECT 275.940 1.400 276.780 1279.600 ;
    RECT 277.060 1.400 277.900 1279.600 ;
    RECT 278.180 1.400 279.020 1279.600 ;
    RECT 279.300 1.400 280.140 1279.600 ;
    RECT 280.420 1.400 281.260 1279.600 ;
    RECT 281.540 1.400 282.380 1279.600 ;
    RECT 282.660 1.400 283.500 1279.600 ;
    RECT 283.780 1.400 284.620 1279.600 ;
    RECT 284.900 1.400 285.740 1279.600 ;
    RECT 286.020 1.400 286.860 1279.600 ;
    RECT 287.140 1.400 287.980 1279.600 ;
    RECT 288.260 1.400 289.100 1279.600 ;
    RECT 289.380 1.400 290.220 1279.600 ;
    RECT 290.500 1.400 291.340 1279.600 ;
    RECT 291.620 1.400 292.460 1279.600 ;
    RECT 292.740 1.400 293.580 1279.600 ;
    RECT 293.860 1.400 294.700 1279.600 ;
    RECT 294.980 1.400 295.820 1279.600 ;
    RECT 296.100 1.400 296.940 1279.600 ;
    RECT 297.220 1.400 298.060 1279.600 ;
    RECT 298.340 1.400 299.180 1279.600 ;
    RECT 299.460 1.400 300.300 1279.600 ;
    RECT 300.580 1.400 301.420 1279.600 ;
    RECT 301.700 1.400 302.540 1279.600 ;
    RECT 302.820 1.400 303.660 1279.600 ;
    RECT 303.940 1.400 304.780 1279.600 ;
    RECT 305.060 1.400 305.900 1279.600 ;
    RECT 306.180 1.400 307.020 1279.600 ;
    RECT 307.300 1.400 308.140 1279.600 ;
    RECT 308.420 1.400 309.260 1279.600 ;
    RECT 309.540 1.400 310.380 1279.600 ;
    RECT 310.660 1.400 311.500 1279.600 ;
    RECT 311.780 1.400 312.620 1279.600 ;
    RECT 312.900 1.400 313.740 1279.600 ;
    RECT 314.020 1.400 314.860 1279.600 ;
    RECT 315.140 1.400 315.980 1279.600 ;
    RECT 316.260 1.400 317.100 1279.600 ;
    RECT 317.380 1.400 318.220 1279.600 ;
    RECT 318.500 1.400 319.340 1279.600 ;
    RECT 319.620 1.400 320.460 1279.600 ;
    RECT 320.740 1.400 321.580 1279.600 ;
    RECT 321.860 1.400 322.700 1279.600 ;
    RECT 322.980 1.400 323.820 1279.600 ;
    RECT 324.100 1.400 324.940 1279.600 ;
    RECT 325.220 1.400 326.060 1279.600 ;
    RECT 326.340 1.400 327.180 1279.600 ;
    RECT 327.460 1.400 328.300 1279.600 ;
    RECT 328.580 1.400 329.420 1279.600 ;
    RECT 329.700 1.400 330.540 1279.600 ;
    RECT 330.820 1.400 331.660 1279.600 ;
    RECT 331.940 1.400 332.780 1279.600 ;
    RECT 333.060 1.400 333.900 1279.600 ;
    RECT 334.180 1.400 335.020 1279.600 ;
    RECT 335.300 1.400 336.140 1279.600 ;
    RECT 336.420 1.400 337.260 1279.600 ;
    RECT 337.540 1.400 338.380 1279.600 ;
    RECT 338.660 1.400 339.500 1279.600 ;
    RECT 339.780 1.400 340.620 1279.600 ;
    RECT 340.900 1.400 341.740 1279.600 ;
    RECT 342.020 1.400 342.860 1279.600 ;
    RECT 343.140 1.400 343.980 1279.600 ;
    RECT 344.260 1.400 345.100 1279.600 ;
    RECT 345.380 1.400 346.220 1279.600 ;
    RECT 346.500 1.400 347.340 1279.600 ;
    RECT 347.620 1.400 348.460 1279.600 ;
    RECT 348.740 1.400 349.580 1279.600 ;
    RECT 349.860 1.400 350.700 1279.600 ;
    RECT 350.980 1.400 351.820 1279.600 ;
    RECT 352.100 1.400 352.940 1279.600 ;
    RECT 353.220 1.400 354.060 1279.600 ;
    RECT 354.340 1.400 355.180 1279.600 ;
    RECT 355.460 1.400 356.300 1279.600 ;
    RECT 356.580 1.400 357.420 1279.600 ;
    RECT 357.700 1.400 358.540 1279.600 ;
    RECT 358.820 1.400 359.660 1279.600 ;
    RECT 359.940 1.400 360.780 1279.600 ;
    RECT 361.060 1.400 361.900 1279.600 ;
    RECT 362.180 1.400 363.020 1279.600 ;
    RECT 363.300 1.400 364.140 1279.600 ;
    RECT 364.420 1.400 365.260 1279.600 ;
    RECT 365.540 1.400 366.380 1279.600 ;
    RECT 366.660 1.400 367.500 1279.600 ;
    RECT 367.780 1.400 368.620 1279.600 ;
    RECT 368.900 1.400 369.740 1279.600 ;
    RECT 370.020 1.400 370.860 1279.600 ;
    RECT 371.140 1.400 371.980 1279.600 ;
    RECT 372.260 1.400 373.100 1279.600 ;
    RECT 373.380 1.400 374.220 1279.600 ;
    RECT 374.500 1.400 375.340 1279.600 ;
    RECT 375.620 1.400 376.460 1279.600 ;
    RECT 376.740 1.400 377.580 1279.600 ;
    RECT 377.860 1.400 378.700 1279.600 ;
    RECT 378.980 1.400 379.820 1279.600 ;
    RECT 380.100 1.400 380.940 1279.600 ;
    RECT 381.220 1.400 382.060 1279.600 ;
    RECT 382.340 1.400 383.180 1279.600 ;
    RECT 383.460 1.400 384.300 1279.600 ;
    RECT 384.580 1.400 385.420 1279.600 ;
    RECT 385.700 1.400 386.540 1279.600 ;
    RECT 386.820 1.400 387.660 1279.600 ;
    RECT 387.940 1.400 388.780 1279.600 ;
    RECT 389.060 1.400 389.900 1279.600 ;
    RECT 390.180 1.400 391.020 1279.600 ;
    RECT 391.300 1.400 392.140 1279.600 ;
    RECT 392.420 1.400 393.260 1279.600 ;
    RECT 393.540 1.400 394.380 1279.600 ;
    RECT 394.660 1.400 395.500 1279.600 ;
    RECT 395.780 1.400 396.620 1279.600 ;
    RECT 396.900 1.400 397.740 1279.600 ;
    RECT 398.020 1.400 398.860 1279.600 ;
    RECT 399.140 1.400 399.980 1279.600 ;
    RECT 400.260 1.400 401.100 1279.600 ;
    RECT 401.380 1.400 402.220 1279.600 ;
    RECT 402.500 1.400 403.340 1279.600 ;
    RECT 403.620 1.400 404.460 1279.600 ;
    RECT 404.740 1.400 405.580 1279.600 ;
    RECT 405.860 1.400 406.700 1279.600 ;
    RECT 406.980 1.400 407.820 1279.600 ;
    RECT 408.100 1.400 408.940 1279.600 ;
    RECT 409.220 1.400 410.060 1279.600 ;
    RECT 410.340 1.400 411.180 1279.600 ;
    RECT 411.460 1.400 412.300 1279.600 ;
    RECT 412.580 1.400 413.420 1279.600 ;
    RECT 413.700 1.400 414.540 1279.600 ;
    RECT 414.820 1.400 415.660 1279.600 ;
    RECT 415.940 1.400 416.780 1279.600 ;
    RECT 417.060 1.400 417.900 1279.600 ;
    RECT 418.180 1.400 419.020 1279.600 ;
    RECT 419.300 1.400 420.140 1279.600 ;
    RECT 420.420 1.400 421.260 1279.600 ;
    RECT 421.540 1.400 422.380 1279.600 ;
    RECT 422.660 1.400 423.500 1279.600 ;
    RECT 423.780 1.400 424.620 1279.600 ;
    RECT 424.900 1.400 425.740 1279.600 ;
    RECT 426.020 1.400 426.860 1279.600 ;
    RECT 427.140 1.400 427.980 1279.600 ;
    RECT 428.260 1.400 429.100 1279.600 ;
    RECT 429.380 1.400 430.220 1279.600 ;
    RECT 430.500 1.400 431.340 1279.600 ;
    RECT 431.620 1.400 432.460 1279.600 ;
    RECT 432.740 1.400 433.580 1279.600 ;
    RECT 433.860 1.400 434.700 1279.600 ;
    RECT 434.980 1.400 435.820 1279.600 ;
    RECT 436.100 1.400 436.940 1279.600 ;
    RECT 437.220 1.400 438.060 1279.600 ;
    RECT 438.340 1.400 439.180 1279.600 ;
    RECT 439.460 1.400 440.300 1279.600 ;
    RECT 440.580 1.400 441.420 1279.600 ;
    RECT 441.700 1.400 442.540 1279.600 ;
    RECT 442.820 1.400 443.660 1279.600 ;
    RECT 443.940 1.400 444.780 1279.600 ;
    RECT 445.060 1.400 445.900 1279.600 ;
    RECT 446.180 1.400 447.020 1279.600 ;
    RECT 447.300 1.400 448.140 1279.600 ;
    RECT 448.420 1.400 449.260 1279.600 ;
    RECT 449.540 1.400 450.380 1279.600 ;
    RECT 450.660 1.400 451.500 1279.600 ;
    RECT 451.780 1.400 452.620 1279.600 ;
    RECT 452.900 1.400 453.740 1279.600 ;
    RECT 454.020 1.400 454.860 1279.600 ;
    RECT 455.140 1.400 455.980 1279.600 ;
    RECT 456.260 1.400 457.100 1279.600 ;
    RECT 457.380 1.400 458.220 1279.600 ;
    RECT 458.500 1.400 459.340 1279.600 ;
    RECT 459.620 1.400 460.460 1279.600 ;
    RECT 460.740 1.400 461.580 1279.600 ;
    RECT 461.860 1.400 462.700 1279.600 ;
    RECT 462.980 1.400 463.820 1279.600 ;
    RECT 464.100 1.400 464.940 1279.600 ;
    RECT 465.220 1.400 466.060 1279.600 ;
    RECT 466.340 1.400 467.180 1279.600 ;
    RECT 467.460 1.400 468.300 1279.600 ;
    RECT 468.580 1.400 469.420 1279.600 ;
    RECT 469.700 1.400 470.540 1279.600 ;
    RECT 470.820 1.400 471.660 1279.600 ;
    RECT 471.940 1.400 472.780 1279.600 ;
    RECT 473.060 1.400 473.900 1279.600 ;
    RECT 474.180 1.400 475.020 1279.600 ;
    RECT 475.300 1.400 476.140 1279.600 ;
    RECT 476.420 1.400 477.260 1279.600 ;
    RECT 477.540 1.400 478.380 1279.600 ;
    RECT 478.660 1.400 479.500 1279.600 ;
    RECT 479.780 1.400 480.620 1279.600 ;
    RECT 480.900 1.400 481.740 1279.600 ;
    RECT 482.020 1.400 482.860 1279.600 ;
    RECT 483.140 1.400 483.980 1279.600 ;
    RECT 484.260 1.400 485.100 1279.600 ;
    RECT 485.380 1.400 486.220 1279.600 ;
    RECT 486.500 1.400 487.340 1279.600 ;
    RECT 487.620 1.400 488.460 1279.600 ;
    RECT 488.740 1.400 489.580 1279.600 ;
    RECT 489.860 1.400 490.700 1279.600 ;
    RECT 490.980 1.400 491.820 1279.600 ;
    RECT 492.100 1.400 492.940 1279.600 ;
    RECT 493.220 1.400 494.060 1279.600 ;
    RECT 494.340 1.400 495.180 1279.600 ;
    RECT 495.460 1.400 496.300 1279.600 ;
    RECT 496.580 1.400 497.420 1279.600 ;
    RECT 497.700 1.400 498.540 1279.600 ;
    RECT 498.820 1.400 499.660 1279.600 ;
    RECT 499.940 1.400 500.780 1279.600 ;
    RECT 501.060 1.400 501.900 1279.600 ;
    RECT 502.180 1.400 503.020 1279.600 ;
    RECT 503.300 1.400 504.140 1279.600 ;
    RECT 504.420 1.400 505.260 1279.600 ;
    RECT 505.540 1.400 506.380 1279.600 ;
    RECT 506.660 1.400 507.500 1279.600 ;
    RECT 507.780 1.400 508.620 1279.600 ;
    RECT 508.900 1.400 509.740 1279.600 ;
    RECT 510.020 1.400 510.860 1279.600 ;
    RECT 511.140 1.400 511.980 1279.600 ;
    RECT 512.260 1.400 513.100 1279.600 ;
    RECT 513.380 1.400 514.220 1279.600 ;
    RECT 514.500 1.400 515.340 1279.600 ;
    RECT 515.620 1.400 516.460 1279.600 ;
    RECT 516.740 1.400 517.580 1279.600 ;
    RECT 517.860 1.400 518.700 1279.600 ;
    RECT 518.980 1.400 519.820 1279.600 ;
    RECT 520.100 1.400 520.940 1279.600 ;
    RECT 521.220 1.400 522.060 1279.600 ;
    RECT 522.340 1.400 523.180 1279.600 ;
    RECT 523.460 1.400 524.300 1279.600 ;
    RECT 524.580 1.400 525.420 1279.600 ;
    RECT 525.700 1.400 526.540 1279.600 ;
    RECT 526.820 1.400 527.660 1279.600 ;
    RECT 527.940 1.400 528.780 1279.600 ;
    RECT 529.060 1.400 529.900 1279.600 ;
    RECT 530.180 1.400 531.020 1279.600 ;
    RECT 531.300 1.400 532.140 1279.600 ;
    RECT 532.420 1.400 533.260 1279.600 ;
    RECT 533.540 1.400 534.380 1279.600 ;
    RECT 534.660 1.400 535.500 1279.600 ;
    RECT 535.780 1.400 536.620 1279.600 ;
    RECT 536.900 1.400 537.740 1279.600 ;
    RECT 538.020 1.400 538.860 1279.600 ;
    RECT 539.140 1.400 539.980 1279.600 ;
    RECT 540.260 1.400 541.100 1279.600 ;
    RECT 541.380 1.400 542.220 1279.600 ;
    RECT 542.500 1.400 543.340 1279.600 ;
    RECT 543.620 1.400 544.460 1279.600 ;
    RECT 544.740 1.400 545.580 1279.600 ;
    RECT 545.860 1.400 546.700 1279.600 ;
    RECT 546.980 1.400 547.820 1279.600 ;
    RECT 548.100 1.400 548.940 1279.600 ;
    RECT 549.220 1.400 550.060 1279.600 ;
    RECT 550.340 1.400 551.180 1279.600 ;
    RECT 551.460 1.400 552.300 1279.600 ;
    RECT 552.580 1.400 553.420 1279.600 ;
    RECT 553.700 1.400 554.540 1279.600 ;
    RECT 554.820 1.400 555.660 1279.600 ;
    RECT 555.940 1.400 556.780 1279.600 ;
    RECT 557.060 1.400 557.900 1279.600 ;
    RECT 558.180 1.400 559.020 1279.600 ;
    RECT 559.300 1.400 560.140 1279.600 ;
    RECT 560.420 1.400 561.260 1279.600 ;
    RECT 561.540 1.400 562.380 1279.600 ;
    RECT 562.660 1.400 563.500 1279.600 ;
    RECT 563.780 1.400 564.620 1279.600 ;
    RECT 564.900 1.400 565.740 1279.600 ;
    RECT 566.020 1.400 566.860 1279.600 ;
    RECT 567.140 1.400 567.980 1279.600 ;
    RECT 568.260 1.400 569.100 1279.600 ;
    RECT 569.380 1.400 570.220 1279.600 ;
    RECT 570.500 1.400 571.340 1279.600 ;
    RECT 571.620 1.400 572.460 1279.600 ;
    RECT 572.740 1.400 573.580 1279.600 ;
    RECT 573.860 1.400 574.700 1279.600 ;
    RECT 574.980 1.400 575.820 1279.600 ;
    RECT 576.100 1.400 576.940 1279.600 ;
    RECT 577.220 1.400 578.060 1279.600 ;
    RECT 578.340 1.400 579.180 1279.600 ;
    RECT 579.460 1.400 580.300 1279.600 ;
    RECT 580.580 1.400 581.420 1279.600 ;
    RECT 581.700 1.400 582.540 1279.600 ;
    RECT 582.820 1.400 583.660 1279.600 ;
    RECT 583.940 1.400 584.780 1279.600 ;
    RECT 585.060 1.400 585.900 1279.600 ;
    RECT 586.180 1.400 587.020 1279.600 ;
    RECT 587.300 1.400 588.140 1279.600 ;
    RECT 588.420 1.400 589.260 1279.600 ;
    RECT 589.540 1.400 590.380 1279.600 ;
    RECT 590.660 1.400 591.500 1279.600 ;
    RECT 591.780 1.400 592.620 1279.600 ;
    RECT 592.900 1.400 593.740 1279.600 ;
    RECT 594.020 1.400 594.860 1279.600 ;
    RECT 595.140 1.400 595.980 1279.600 ;
    RECT 596.260 1.400 597.100 1279.600 ;
    RECT 597.380 1.400 598.220 1279.600 ;
    RECT 598.500 1.400 599.340 1279.600 ;
    RECT 599.620 1.400 600.460 1279.600 ;
    RECT 600.740 1.400 601.580 1279.600 ;
    RECT 601.860 1.400 602.700 1279.600 ;
    RECT 602.980 1.400 603.820 1279.600 ;
    RECT 604.100 1.400 604.940 1279.600 ;
    RECT 605.220 1.400 606.060 1279.600 ;
    RECT 606.340 1.400 607.180 1279.600 ;
    RECT 607.460 1.400 608.300 1279.600 ;
    RECT 608.580 1.400 609.420 1279.600 ;
    RECT 609.700 1.400 610.540 1279.600 ;
    RECT 610.820 1.400 611.660 1279.600 ;
    RECT 611.940 1.400 612.780 1279.600 ;
    RECT 613.060 1.400 613.900 1279.600 ;
    RECT 614.180 1.400 615.020 1279.600 ;
    RECT 615.300 1.400 616.140 1279.600 ;
    RECT 616.420 1.400 617.260 1279.600 ;
    RECT 617.540 1.400 618.380 1279.600 ;
    RECT 618.660 1.400 619.500 1279.600 ;
    RECT 619.780 1.400 620.620 1279.600 ;
    RECT 620.900 1.400 621.740 1279.600 ;
    RECT 622.020 1.400 622.860 1279.600 ;
    RECT 623.140 1.400 623.980 1279.600 ;
    RECT 624.260 1.400 625.100 1279.600 ;
    RECT 625.380 1.400 626.220 1279.600 ;
    RECT 626.500 1.400 627.340 1279.600 ;
    RECT 627.620 1.400 628.460 1279.600 ;
    RECT 628.740 1.400 629.580 1279.600 ;
    RECT 629.860 1.400 630.700 1279.600 ;
    RECT 630.980 1.400 631.820 1279.600 ;
    RECT 632.100 1.400 632.940 1279.600 ;
    RECT 633.220 1.400 634.060 1279.600 ;
    RECT 634.340 1.400 635.180 1279.600 ;
    RECT 635.460 1.400 636.300 1279.600 ;
    RECT 636.580 1.400 637.420 1279.600 ;
    RECT 637.700 1.400 638.540 1279.600 ;
    RECT 638.820 1.400 639.660 1279.600 ;
    RECT 639.940 1.400 640.780 1279.600 ;
    RECT 641.060 1.400 641.900 1279.600 ;
    RECT 642.180 1.400 643.020 1279.600 ;
    RECT 643.300 1.400 644.140 1279.600 ;
    RECT 644.420 1.400 645.260 1279.600 ;
    RECT 645.540 1.400 646.380 1279.600 ;
    RECT 646.660 1.400 647.500 1279.600 ;
    RECT 647.780 1.400 648.620 1279.600 ;
    RECT 648.900 1.400 649.740 1279.600 ;
    RECT 650.020 1.400 650.860 1279.600 ;
    RECT 651.140 1.400 651.980 1279.600 ;
    RECT 652.260 1.400 653.100 1279.600 ;
    RECT 653.380 1.400 654.220 1279.600 ;
    RECT 654.500 1.400 655.340 1279.600 ;
    RECT 655.620 1.400 656.460 1279.600 ;
    RECT 656.740 1.400 657.580 1279.600 ;
    RECT 657.860 1.400 658.700 1279.600 ;
    RECT 658.980 1.400 659.820 1279.600 ;
    RECT 660.100 1.400 660.940 1279.600 ;
    RECT 661.220 1.400 662.060 1279.600 ;
    RECT 662.340 1.400 663.180 1279.600 ;
    RECT 663.460 1.400 664.300 1279.600 ;
    RECT 664.580 1.400 665.420 1279.600 ;
    RECT 665.700 1.400 666.540 1279.600 ;
    RECT 666.820 1.400 667.660 1279.600 ;
    RECT 667.940 1.400 668.780 1279.600 ;
    RECT 669.060 1.400 669.900 1279.600 ;
    RECT 670.180 1.400 671.020 1279.600 ;
    RECT 671.300 1.400 672.140 1279.600 ;
    RECT 672.420 1.400 673.260 1279.600 ;
    RECT 673.540 1.400 674.380 1279.600 ;
    RECT 674.660 1.400 675.500 1279.600 ;
    RECT 675.780 1.400 676.620 1279.600 ;
    RECT 676.900 1.400 677.740 1279.600 ;
    RECT 678.020 1.400 678.860 1279.600 ;
    RECT 679.140 1.400 679.980 1279.600 ;
    RECT 680.260 1.400 681.100 1279.600 ;
    RECT 681.380 1.400 682.220 1279.600 ;
    RECT 682.500 1.400 683.340 1279.600 ;
    RECT 683.620 1.400 684.460 1279.600 ;
    RECT 684.740 1.400 685.580 1279.600 ;
    RECT 685.860 1.400 686.700 1279.600 ;
    RECT 686.980 1.400 687.820 1279.600 ;
    RECT 688.100 1.400 688.940 1279.600 ;
    RECT 689.220 1.400 690.060 1279.600 ;
    RECT 690.340 1.400 691.180 1279.600 ;
    RECT 691.460 1.400 692.300 1279.600 ;
    RECT 692.580 1.400 693.420 1279.600 ;
    RECT 693.700 1.400 694.540 1279.600 ;
    RECT 694.820 1.400 695.660 1279.600 ;
    RECT 695.940 1.400 696.780 1279.600 ;
    RECT 697.060 1.400 697.900 1279.600 ;
    RECT 698.180 1.400 699.020 1279.600 ;
    RECT 699.300 1.400 700.140 1279.600 ;
    RECT 700.420 1.400 701.260 1279.600 ;
    RECT 701.540 1.400 702.380 1279.600 ;
    RECT 702.660 1.400 703.500 1279.600 ;
    RECT 703.780 1.400 704.620 1279.600 ;
    RECT 704.900 1.400 705.740 1279.600 ;
    RECT 706.020 1.400 706.860 1279.600 ;
    RECT 707.140 1.400 707.980 1279.600 ;
    RECT 708.260 1.400 709.100 1279.600 ;
    RECT 709.380 1.400 710.220 1279.600 ;
    RECT 710.500 1.400 711.340 1279.600 ;
    RECT 711.620 1.400 712.460 1279.600 ;
    RECT 712.740 1.400 713.580 1279.600 ;
    RECT 713.860 1.400 714.700 1279.600 ;
    RECT 714.980 1.400 715.820 1279.600 ;
    RECT 716.100 1.400 716.940 1279.600 ;
    RECT 717.220 1.400 718.060 1279.600 ;
    RECT 718.340 1.400 719.180 1279.600 ;
    RECT 719.460 1.400 720.300 1279.600 ;
    RECT 720.580 1.400 721.420 1279.600 ;
    RECT 721.700 1.400 722.540 1279.600 ;
    RECT 722.820 1.400 723.660 1279.600 ;
    RECT 723.940 1.400 724.780 1279.600 ;
    RECT 725.060 1.400 725.900 1279.600 ;
    RECT 726.180 1.400 727.020 1279.600 ;
    RECT 727.300 1.400 728.140 1279.600 ;
    RECT 728.420 1.400 729.260 1279.600 ;
    RECT 729.540 1.400 730.380 1279.600 ;
    RECT 730.660 1.400 731.500 1279.600 ;
    RECT 731.780 1.400 732.620 1279.600 ;
    RECT 732.900 1.400 733.740 1279.600 ;
    RECT 734.020 1.400 734.860 1279.600 ;
    RECT 735.140 1.400 735.980 1279.600 ;
    RECT 736.260 1.400 737.100 1279.600 ;
    RECT 737.380 1.400 738.220 1279.600 ;
    RECT 738.500 1.400 739.340 1279.600 ;
    RECT 739.620 1.400 740.460 1279.600 ;
    RECT 740.740 1.400 741.580 1279.600 ;
    RECT 741.860 1.400 742.700 1279.600 ;
    RECT 742.980 1.400 743.820 1279.600 ;
    RECT 744.100 1.400 744.940 1279.600 ;
    RECT 745.220 1.400 746.060 1279.600 ;
    RECT 746.340 1.400 747.180 1279.600 ;
    RECT 747.460 1.400 748.300 1279.600 ;
    RECT 748.580 1.400 749.420 1279.600 ;
    RECT 749.700 1.400 750.540 1279.600 ;
    RECT 750.820 1.400 751.660 1279.600 ;
    RECT 751.940 1.400 752.780 1279.600 ;
    RECT 753.060 1.400 753.900 1279.600 ;
    RECT 754.180 1.400 755.020 1279.600 ;
    RECT 755.300 1.400 756.140 1279.600 ;
    RECT 756.420 1.400 757.260 1279.600 ;
    RECT 757.540 1.400 758.380 1279.600 ;
    RECT 758.660 1.400 759.500 1279.600 ;
    RECT 759.780 1.400 760.620 1279.600 ;
    RECT 760.900 1.400 761.740 1279.600 ;
    RECT 762.020 1.400 762.860 1279.600 ;
    RECT 763.140 1.400 763.980 1279.600 ;
    RECT 764.260 1.400 765.100 1279.600 ;
    RECT 765.380 1.400 766.220 1279.600 ;
    RECT 766.500 1.400 767.340 1279.600 ;
    RECT 767.620 1.400 768.460 1279.600 ;
    RECT 768.740 1.400 769.580 1279.600 ;
    RECT 769.860 1.400 770.700 1279.600 ;
    RECT 770.980 1.400 771.820 1279.600 ;
    RECT 772.100 1.400 772.940 1279.600 ;
    RECT 773.220 1.400 774.060 1279.600 ;
    RECT 774.340 1.400 775.180 1279.600 ;
    RECT 775.460 1.400 776.300 1279.600 ;
    RECT 776.580 1.400 777.420 1279.600 ;
    RECT 777.700 1.400 778.540 1279.600 ;
    RECT 778.820 1.400 779.660 1279.600 ;
    RECT 779.940 1.400 780.780 1279.600 ;
    RECT 781.060 1.400 781.900 1279.600 ;
    RECT 782.180 1.400 783.020 1279.600 ;
    RECT 783.300 1.400 784.140 1279.600 ;
    RECT 784.420 1.400 785.260 1279.600 ;
    RECT 785.540 1.400 786.380 1279.600 ;
    RECT 786.660 1.400 787.500 1279.600 ;
    RECT 787.780 1.400 788.620 1279.600 ;
    RECT 788.900 1.400 789.740 1279.600 ;
    RECT 790.020 1.400 790.860 1279.600 ;
    RECT 791.140 1.400 791.980 1279.600 ;
    RECT 792.260 1.400 793.100 1279.600 ;
    RECT 793.380 1.400 794.220 1279.600 ;
    RECT 794.500 1.400 795.340 1279.600 ;
    RECT 795.620 1.400 796.460 1279.600 ;
    RECT 796.740 1.400 797.580 1279.600 ;
    RECT 797.860 1.400 798.700 1279.600 ;
    RECT 798.980 1.400 799.820 1279.600 ;
    RECT 800.100 1.400 800.940 1279.600 ;
    RECT 801.220 1.400 802.060 1279.600 ;
    RECT 802.340 1.400 803.180 1279.600 ;
    RECT 803.460 1.400 804.300 1279.600 ;
    RECT 804.580 1.400 805.420 1279.600 ;
    RECT 805.700 1.400 806.540 1279.600 ;
    RECT 806.820 1.400 807.660 1279.600 ;
    RECT 807.940 1.400 808.780 1279.600 ;
    RECT 809.060 1.400 809.900 1279.600 ;
    RECT 810.180 1.400 811.020 1279.600 ;
    RECT 811.300 1.400 812.140 1279.600 ;
    RECT 812.420 1.400 813.260 1279.600 ;
    RECT 813.540 1.400 814.380 1279.600 ;
    RECT 814.660 1.400 815.500 1279.600 ;
    RECT 815.780 1.400 816.620 1279.600 ;
    RECT 816.900 1.400 817.740 1279.600 ;
    RECT 818.020 1.400 818.860 1279.600 ;
    RECT 819.140 1.400 819.980 1279.600 ;
    RECT 820.260 1.400 821.100 1279.600 ;
    RECT 821.380 1.400 822.220 1279.600 ;
    RECT 822.500 1.400 823.340 1279.600 ;
    RECT 823.620 1.400 824.460 1279.600 ;
    RECT 824.740 1.400 825.580 1279.600 ;
    RECT 825.860 1.400 826.700 1279.600 ;
    RECT 826.980 1.400 827.820 1279.600 ;
    RECT 828.100 1.400 828.940 1279.600 ;
    RECT 829.220 1.400 830.060 1279.600 ;
    RECT 830.340 1.400 831.180 1279.600 ;
    RECT 831.460 1.400 832.300 1279.600 ;
    RECT 832.580 1.400 833.420 1279.600 ;
    RECT 833.700 1.400 834.540 1279.600 ;
    RECT 834.820 1.400 835.660 1279.600 ;
    RECT 835.940 1.400 836.780 1279.600 ;
    RECT 837.060 1.400 837.900 1279.600 ;
    RECT 838.180 1.400 839.020 1279.600 ;
    RECT 839.300 1.400 840.140 1279.600 ;
    RECT 840.420 1.400 841.260 1279.600 ;
    RECT 841.540 1.400 842.380 1279.600 ;
    RECT 842.660 1.400 843.500 1279.600 ;
    RECT 843.780 1.400 844.620 1279.600 ;
    RECT 844.900 1.400 845.740 1279.600 ;
    RECT 846.020 1.400 846.860 1279.600 ;
    RECT 847.140 1.400 847.980 1279.600 ;
    RECT 848.260 1.400 849.100 1279.600 ;
    RECT 849.380 1.400 850.220 1279.600 ;
    RECT 850.500 1.400 851.340 1279.600 ;
    RECT 851.620 1.400 852.460 1279.600 ;
    RECT 852.740 1.400 853.580 1279.600 ;
    RECT 853.860 1.400 854.700 1279.600 ;
    RECT 854.980 1.400 855.820 1279.600 ;
    RECT 856.100 1.400 856.940 1279.600 ;
    RECT 857.220 1.400 858.060 1279.600 ;
    RECT 858.340 1.400 859.180 1279.600 ;
    RECT 859.460 1.400 860.300 1279.600 ;
    RECT 860.580 1.400 861.420 1279.600 ;
    RECT 861.700 1.400 862.540 1279.600 ;
    RECT 862.820 1.400 863.660 1279.600 ;
    RECT 863.940 1.400 864.780 1279.600 ;
    RECT 865.060 1.400 865.900 1279.600 ;
    RECT 866.180 1.400 867.020 1279.600 ;
    RECT 867.300 1.400 868.140 1279.600 ;
    RECT 868.420 1.400 869.260 1279.600 ;
    RECT 869.540 1.400 870.380 1279.600 ;
    RECT 870.660 1.400 871.500 1279.600 ;
    RECT 871.780 1.400 872.620 1279.600 ;
    RECT 872.900 1.400 873.740 1279.600 ;
    RECT 874.020 1.400 874.860 1279.600 ;
    RECT 875.140 1.400 875.980 1279.600 ;
    RECT 876.260 1.400 877.100 1279.600 ;
    RECT 877.380 1.400 878.220 1279.600 ;
    RECT 878.500 1.400 879.340 1279.600 ;
    RECT 879.620 1.400 880.460 1279.600 ;
    RECT 880.740 1.400 881.580 1279.600 ;
    RECT 881.860 1.400 882.700 1279.600 ;
    RECT 882.980 1.400 883.820 1279.600 ;
    RECT 884.100 1.400 884.940 1279.600 ;
    RECT 885.220 1.400 886.060 1279.600 ;
    RECT 886.340 1.400 887.180 1279.600 ;
    RECT 887.460 1.400 888.300 1279.600 ;
    RECT 888.580 1.400 889.420 1279.600 ;
    RECT 889.700 1.400 890.540 1279.600 ;
    RECT 890.820 1.400 891.660 1279.600 ;
    RECT 891.940 1.400 892.780 1279.600 ;
    RECT 893.060 1.400 893.900 1279.600 ;
    RECT 894.180 1.400 895.020 1279.600 ;
    RECT 895.300 1.400 896.140 1279.600 ;
    RECT 896.420 1.400 897.260 1279.600 ;
    RECT 897.540 1.400 898.380 1279.600 ;
    RECT 898.660 1.400 899.500 1279.600 ;
    RECT 899.780 1.400 900.620 1279.600 ;
    RECT 900.900 1.400 901.740 1279.600 ;
    RECT 902.020 1.400 902.860 1279.600 ;
    RECT 903.140 1.400 903.980 1279.600 ;
    RECT 904.260 1.400 905.100 1279.600 ;
    RECT 905.380 1.400 906.220 1279.600 ;
    RECT 906.500 1.400 907.340 1279.600 ;
    RECT 907.620 1.400 908.460 1279.600 ;
    RECT 908.740 1.400 909.580 1279.600 ;
    RECT 909.860 1.400 910.700 1279.600 ;
    RECT 910.980 1.400 911.820 1279.600 ;
    RECT 912.100 1.400 912.940 1279.600 ;
    RECT 913.220 1.400 914.060 1279.600 ;
    RECT 914.340 1.400 915.180 1279.600 ;
    RECT 915.460 1.400 916.300 1279.600 ;
    RECT 916.580 1.400 917.420 1279.600 ;
    RECT 917.700 1.400 918.540 1279.600 ;
    RECT 918.820 1.400 919.660 1279.600 ;
    RECT 919.940 1.400 920.780 1279.600 ;
    RECT 921.060 1.400 921.900 1279.600 ;
    RECT 922.180 1.400 923.020 1279.600 ;
    RECT 923.300 1.400 924.140 1279.600 ;
    RECT 924.420 1.400 925.260 1279.600 ;
    RECT 925.540 1.400 926.380 1279.600 ;
    RECT 926.660 1.400 927.500 1279.600 ;
    RECT 927.780 1.400 928.620 1279.600 ;
    RECT 928.900 1.400 929.740 1279.600 ;
    RECT 930.020 1.400 930.860 1279.600 ;
    RECT 931.140 1.400 931.980 1279.600 ;
    RECT 932.260 1.400 933.100 1279.600 ;
    RECT 933.380 1.400 934.220 1279.600 ;
    RECT 934.500 1.400 935.340 1279.600 ;
    RECT 935.620 1.400 936.460 1279.600 ;
    RECT 936.740 1.400 937.580 1279.600 ;
    RECT 937.860 1.400 938.700 1279.600 ;
    RECT 938.980 1.400 939.820 1279.600 ;
    RECT 940.100 1.400 940.940 1279.600 ;
    RECT 941.220 1.400 942.060 1279.600 ;
    RECT 942.340 1.400 943.180 1279.600 ;
    RECT 943.460 1.400 944.300 1279.600 ;
    RECT 944.580 1.400 945.420 1279.600 ;
    RECT 945.700 1.400 946.540 1279.600 ;
    RECT 946.820 1.400 947.660 1279.600 ;
    RECT 947.940 1.400 948.780 1279.600 ;
    RECT 949.060 1.400 949.900 1279.600 ;
    RECT 950.180 1.400 951.020 1279.600 ;
    RECT 951.300 1.400 952.140 1279.600 ;
    RECT 952.420 1.400 953.260 1279.600 ;
    RECT 953.540 1.400 954.380 1279.600 ;
    RECT 954.660 1.400 955.500 1279.600 ;
    RECT 955.780 1.400 956.620 1279.600 ;
    RECT 956.900 1.400 957.740 1279.600 ;
    RECT 958.020 1.400 958.860 1279.600 ;
    RECT 959.140 1.400 959.980 1279.600 ;
    RECT 960.260 1.400 961.100 1279.600 ;
    RECT 961.380 1.400 962.220 1279.600 ;
    RECT 962.500 1.400 963.340 1279.600 ;
    RECT 963.620 1.400 964.460 1279.600 ;
    RECT 964.740 1.400 965.580 1279.600 ;
    RECT 965.860 1.400 966.700 1279.600 ;
    RECT 966.980 1.400 967.820 1279.600 ;
    RECT 968.100 1.400 968.940 1279.600 ;
    RECT 969.220 1.400 970.060 1279.600 ;
    RECT 970.340 1.400 971.180 1279.600 ;
    RECT 971.460 1.400 972.300 1279.600 ;
    RECT 972.580 1.400 973.420 1279.600 ;
    RECT 973.700 1.400 974.540 1279.600 ;
    RECT 974.820 1.400 975.660 1279.600 ;
    RECT 975.940 1.400 976.780 1279.600 ;
    RECT 977.060 1.400 977.900 1279.600 ;
    RECT 978.180 1.400 979.020 1279.600 ;
    RECT 979.300 1.400 980.140 1279.600 ;
    RECT 980.420 1.400 981.260 1279.600 ;
    RECT 981.540 1.400 982.380 1279.600 ;
    RECT 982.660 1.400 983.500 1279.600 ;
    RECT 983.780 1.400 984.620 1279.600 ;
    RECT 984.900 1.400 985.740 1279.600 ;
    RECT 986.020 1.400 986.860 1279.600 ;
    RECT 987.140 1.400 987.980 1279.600 ;
    RECT 988.260 1.400 989.100 1279.600 ;
    RECT 989.380 1.400 990.220 1279.600 ;
    RECT 990.500 1.400 991.340 1279.600 ;
    RECT 991.620 1.400 992.460 1279.600 ;
    RECT 992.740 1.400 993.580 1279.600 ;
    RECT 993.860 1.400 994.700 1279.600 ;
    RECT 994.980 1.400 995.820 1279.600 ;
    RECT 996.100 1.400 996.940 1279.600 ;
    RECT 997.220 1.400 998.060 1279.600 ;
    RECT 998.340 1.400 999.180 1279.600 ;
    RECT 999.460 1.400 1000.300 1279.600 ;
    RECT 1000.580 1.400 1001.420 1279.600 ;
    RECT 1001.700 1.400 1002.540 1279.600 ;
    RECT 1002.820 1.400 1003.660 1279.600 ;
    RECT 1003.940 1.400 1004.780 1279.600 ;
    RECT 1005.060 1.400 1005.900 1279.600 ;
    RECT 1006.180 1.400 1007.020 1279.600 ;
    RECT 1007.300 1.400 1008.140 1279.600 ;
    RECT 1008.420 1.400 1009.260 1279.600 ;
    RECT 1009.540 1.400 1010.380 1279.600 ;
    RECT 1010.660 1.400 1011.500 1279.600 ;
    RECT 1011.780 1.400 1012.620 1279.600 ;
    RECT 1012.900 1.400 1013.740 1279.600 ;
    RECT 1014.020 1.400 1014.860 1279.600 ;
    RECT 1015.140 1.400 1015.980 1279.600 ;
    RECT 1016.260 1.400 1017.100 1279.600 ;
    RECT 1017.380 1.400 1018.220 1279.600 ;
    RECT 1018.500 1.400 1019.340 1279.600 ;
    RECT 1019.620 1.400 1020.460 1279.600 ;
    RECT 1020.740 1.400 1021.580 1279.600 ;
    RECT 1021.860 1.400 1022.700 1279.600 ;
    RECT 1022.980 1.400 1023.820 1279.600 ;
    RECT 1024.100 1.400 1024.940 1279.600 ;
    RECT 1025.220 1.400 1026.060 1279.600 ;
    RECT 1026.340 1.400 1027.180 1279.600 ;
    RECT 1027.460 1.400 1028.300 1279.600 ;
    RECT 1028.580 1.400 1029.420 1279.600 ;
    RECT 1029.700 1.400 1030.540 1279.600 ;
    RECT 1030.820 1.400 1031.660 1279.600 ;
    RECT 1031.940 1.400 1032.780 1279.600 ;
    RECT 1033.060 1.400 1033.900 1279.600 ;
    RECT 1034.180 1.400 1035.020 1279.600 ;
    RECT 1035.300 1.400 1036.140 1279.600 ;
    RECT 1036.420 1.400 1037.260 1279.600 ;
    RECT 1037.540 1.400 1038.380 1279.600 ;
    RECT 1038.660 1.400 1039.500 1279.600 ;
    RECT 1039.780 1.400 1040.620 1279.600 ;
    RECT 1040.900 1.400 1041.740 1279.600 ;
    RECT 1042.020 1.400 1042.860 1279.600 ;
    RECT 1043.140 1.400 1043.980 1279.600 ;
    RECT 1044.260 1.400 1045.100 1279.600 ;
    RECT 1045.380 1.400 1046.220 1279.600 ;
    RECT 1046.500 1.400 1047.340 1279.600 ;
    RECT 1047.620 1.400 1048.460 1279.600 ;
    RECT 1048.740 1.400 1049.580 1279.600 ;
    RECT 1049.860 1.400 1050.700 1279.600 ;
    RECT 1050.980 1.400 1051.820 1279.600 ;
    RECT 1052.100 1.400 1052.940 1279.600 ;
    RECT 1053.220 1.400 1054.060 1279.600 ;
    RECT 1054.340 1.400 1055.180 1279.600 ;
    RECT 1055.460 1.400 1056.300 1279.600 ;
    RECT 1056.580 1.400 1057.420 1279.600 ;
    RECT 1057.700 1.400 1058.540 1279.600 ;
    RECT 1058.820 1.400 1059.660 1279.600 ;
    RECT 1059.940 1.400 1060.780 1279.600 ;
    RECT 1061.060 1.400 1061.900 1279.600 ;
    RECT 1062.180 1.400 1063.020 1279.600 ;
    RECT 1063.300 1.400 1064.140 1279.600 ;
    RECT 1064.420 1.400 1065.260 1279.600 ;
    RECT 1065.540 1.400 1066.380 1279.600 ;
    RECT 1066.660 1.400 1067.500 1279.600 ;
    RECT 1067.780 1.400 1068.620 1279.600 ;
    RECT 1068.900 1.400 1069.740 1279.600 ;
    RECT 1070.020 1.400 1070.860 1279.600 ;
    RECT 1071.140 1.400 1071.980 1279.600 ;
    RECT 1072.260 1.400 1073.100 1279.600 ;
    RECT 1073.380 1.400 1074.220 1279.600 ;
    RECT 1074.500 1.400 1075.340 1279.600 ;
    RECT 1075.620 1.400 1076.460 1279.600 ;
    RECT 1076.740 1.400 1077.580 1279.600 ;
    RECT 1077.860 1.400 1078.700 1279.600 ;
    RECT 1078.980 1.400 1079.820 1279.600 ;
    RECT 1080.100 1.400 1080.940 1279.600 ;
    RECT 1081.220 1.400 1082.060 1279.600 ;
    RECT 1082.340 1.400 1083.180 1279.600 ;
    RECT 1083.460 1.400 1084.300 1279.600 ;
    RECT 1084.580 1.400 1085.420 1279.600 ;
    RECT 1085.700 1.400 1086.540 1279.600 ;
    RECT 1086.820 1.400 1087.660 1279.600 ;
    RECT 1087.940 1.400 1088.780 1279.600 ;
    RECT 1089.060 1.400 1089.900 1279.600 ;
    RECT 1090.180 1.400 1091.020 1279.600 ;
    RECT 1091.300 1.400 1092.140 1279.600 ;
    RECT 1092.420 1.400 1093.260 1279.600 ;
    RECT 1093.540 1.400 1094.380 1279.600 ;
    RECT 1094.660 1.400 1095.500 1279.600 ;
    RECT 1095.780 1.400 1096.620 1279.600 ;
    RECT 1096.900 1.400 1097.740 1279.600 ;
    RECT 1098.020 1.400 1098.860 1279.600 ;
    RECT 1099.140 1.400 1099.980 1279.600 ;
    RECT 1100.260 1.400 1101.100 1279.600 ;
    RECT 1101.380 1.400 1102.220 1279.600 ;
    RECT 1102.500 1.400 1103.340 1279.600 ;
    RECT 1103.620 1.400 1104.460 1279.600 ;
    RECT 1104.740 1.400 1105.580 1279.600 ;
    RECT 1105.860 1.400 1106.700 1279.600 ;
    RECT 1106.980 1.400 1107.820 1279.600 ;
    RECT 1108.100 1.400 1108.940 1279.600 ;
    RECT 1109.220 1.400 1110.060 1279.600 ;
    RECT 1110.340 1.400 1111.180 1279.600 ;
    RECT 1111.460 1.400 1112.300 1279.600 ;
    RECT 1112.580 1.400 1113.420 1279.600 ;
    RECT 1113.700 1.400 1114.540 1279.600 ;
    RECT 1114.820 1.400 1115.660 1279.600 ;
    RECT 1115.940 1.400 1116.780 1279.600 ;
    RECT 1117.060 1.400 1117.900 1279.600 ;
    RECT 1118.180 1.400 1119.020 1279.600 ;
    RECT 1119.300 1.400 1120.140 1279.600 ;
    RECT 1120.420 1.400 1121.260 1279.600 ;
    RECT 1121.540 1.400 1122.380 1279.600 ;
    RECT 1122.660 1.400 1123.500 1279.600 ;
    RECT 1123.780 1.400 1124.620 1279.600 ;
    RECT 1124.900 1.400 1125.740 1279.600 ;
    RECT 1126.020 1.400 1126.860 1279.600 ;
    RECT 1127.140 1.400 1127.980 1279.600 ;
    RECT 1128.260 1.400 1129.100 1279.600 ;
    RECT 1129.380 1.400 1130.220 1279.600 ;
    RECT 1130.500 1.400 1131.340 1279.600 ;
    RECT 1131.620 1.400 1132.460 1279.600 ;
    RECT 1132.740 1.400 1133.580 1279.600 ;
    RECT 1133.860 1.400 1134.700 1279.600 ;
    RECT 1134.980 1.400 1135.820 1279.600 ;
    RECT 1136.100 1.400 1136.940 1279.600 ;
    RECT 1137.220 1.400 1138.060 1279.600 ;
    RECT 1138.340 1.400 1139.180 1279.600 ;
    RECT 1139.460 1.400 1140.300 1279.600 ;
    RECT 1140.580 1.400 1141.420 1279.600 ;
    RECT 1141.700 1.400 1142.540 1279.600 ;
    RECT 1142.820 1.400 1143.660 1279.600 ;
    RECT 1143.940 1.400 1144.780 1279.600 ;
    RECT 1145.060 1.400 1145.900 1279.600 ;
    RECT 1146.180 1.400 1147.020 1279.600 ;
    RECT 1147.300 1.400 1148.140 1279.600 ;
    RECT 1148.420 1.400 1149.260 1279.600 ;
    RECT 1149.540 1.400 1150.380 1279.600 ;
    RECT 1150.660 1.400 1151.500 1279.600 ;
    RECT 1151.780 1.400 1152.620 1279.600 ;
    RECT 1152.900 1.400 1153.740 1279.600 ;
    RECT 1154.020 1.400 1154.860 1279.600 ;
    RECT 1155.140 1.400 1155.980 1279.600 ;
    RECT 1156.260 1.400 1157.100 1279.600 ;
    RECT 1157.380 1.400 1158.220 1279.600 ;
    RECT 1158.500 1.400 1159.340 1279.600 ;
    RECT 1159.620 1.400 1160.460 1279.600 ;
    RECT 1160.740 1.400 1161.580 1279.600 ;
    RECT 1161.860 1.400 1162.700 1279.600 ;
    RECT 1162.980 1.400 1163.820 1279.600 ;
    RECT 1164.100 1.400 1164.940 1279.600 ;
    RECT 1165.220 1.400 1166.060 1279.600 ;
    RECT 1166.340 1.400 1167.180 1279.600 ;
    RECT 1167.460 1.400 1168.300 1279.600 ;
    RECT 1168.580 1.400 1169.420 1279.600 ;
    RECT 1169.700 1.400 1170.540 1279.600 ;
    RECT 1170.820 1.400 1171.660 1279.600 ;
    RECT 1171.940 1.400 1172.780 1279.600 ;
    RECT 1173.060 1.400 1173.900 1279.600 ;
    RECT 1174.180 1.400 1175.020 1279.600 ;
    RECT 1175.300 1.400 1176.140 1279.600 ;
    RECT 1176.420 1.400 1177.260 1279.600 ;
    RECT 1177.540 1.400 1178.380 1279.600 ;
    RECT 1178.660 1.400 1179.500 1279.600 ;
    RECT 1179.780 1.400 1180.620 1279.600 ;
    RECT 1180.900 1.400 1181.740 1279.600 ;
    RECT 1182.020 1.400 1182.860 1279.600 ;
    RECT 1183.140 1.400 1183.980 1279.600 ;
    RECT 1184.260 1.400 1185.100 1279.600 ;
    RECT 1185.380 1.400 1186.220 1279.600 ;
    RECT 1186.500 1.400 1187.340 1279.600 ;
    RECT 1187.620 1.400 1188.460 1279.600 ;
    RECT 1188.740 1.400 1189.580 1279.600 ;
    RECT 1189.860 1.400 1190.700 1279.600 ;
    RECT 1190.980 1.400 1191.820 1279.600 ;
    RECT 1192.100 1.400 1192.940 1279.600 ;
    RECT 1193.220 1.400 1194.060 1279.600 ;
    RECT 1194.340 1.400 1195.180 1279.600 ;
    RECT 1195.460 1.400 1196.300 1279.600 ;
    RECT 1196.580 1.400 1197.420 1279.600 ;
    RECT 1197.700 1.400 1198.540 1279.600 ;
    RECT 1198.820 1.400 1199.660 1279.600 ;
    RECT 1199.940 1.400 1200.780 1279.600 ;
    RECT 1201.060 1.400 1201.900 1279.600 ;
    RECT 1202.180 1.400 1203.020 1279.600 ;
    RECT 1203.300 1.400 1204.140 1279.600 ;
    RECT 1204.420 1.400 1205.260 1279.600 ;
    RECT 1205.540 1.400 1206.380 1279.600 ;
    RECT 1206.660 1.400 1207.500 1279.600 ;
    RECT 1207.780 1.400 1208.620 1279.600 ;
    RECT 1208.900 1.400 1209.740 1279.600 ;
    RECT 1210.020 1.400 1210.860 1279.600 ;
    RECT 1211.140 1.400 1211.980 1279.600 ;
    RECT 1212.260 1.400 1213.100 1279.600 ;
    RECT 1213.380 1.400 1214.220 1279.600 ;
    RECT 1214.500 1.400 1215.340 1279.600 ;
    RECT 1215.620 1.400 1216.460 1279.600 ;
    RECT 1216.740 1.400 1217.580 1279.600 ;
    RECT 1217.860 1.400 1218.700 1279.600 ;
    RECT 1218.980 1.400 1219.820 1279.600 ;
    RECT 1220.100 1.400 1220.940 1279.600 ;
    RECT 1221.220 1.400 1222.060 1279.600 ;
    RECT 1222.340 1.400 1223.180 1279.600 ;
    RECT 1223.460 1.400 1224.300 1279.600 ;
    RECT 1224.580 1.400 1225.420 1279.600 ;
    RECT 1225.700 1.400 1226.540 1279.600 ;
    RECT 1226.820 1.400 1227.660 1279.600 ;
    RECT 1227.940 1.400 1228.780 1279.600 ;
    RECT 1229.060 1.400 1229.900 1279.600 ;
    RECT 1230.180 1.400 1231.020 1279.600 ;
    RECT 1231.300 1.400 1232.140 1279.600 ;
    RECT 1232.420 1.400 1233.260 1279.600 ;
    RECT 1233.540 1.400 1234.380 1279.600 ;
    RECT 1234.660 1.400 1235.500 1279.600 ;
    RECT 1235.780 1.400 1236.620 1279.600 ;
    RECT 1236.900 1.400 1237.740 1279.600 ;
    RECT 1238.020 1.400 1238.860 1279.600 ;
    RECT 1239.140 1.400 1239.980 1279.600 ;
    RECT 1240.260 1.400 1241.100 1279.600 ;
    RECT 1241.380 1.400 1242.220 1279.600 ;
    RECT 1242.500 1.400 1243.340 1279.600 ;
    RECT 1243.620 1.400 1244.460 1279.600 ;
    RECT 1244.740 1.400 1245.580 1279.600 ;
    RECT 1245.860 1.400 1246.700 1279.600 ;
    RECT 1246.980 1.400 1247.820 1279.600 ;
    RECT 1248.100 1.400 1248.940 1279.600 ;
    RECT 1249.220 1.400 1250.060 1279.600 ;
    RECT 1250.340 1.400 1251.180 1279.600 ;
    RECT 1251.460 1.400 1252.300 1279.600 ;
    RECT 1252.580 1.400 1253.420 1279.600 ;
    RECT 1253.700 1.400 1254.540 1279.600 ;
    RECT 1254.820 1.400 1255.660 1279.600 ;
    RECT 1255.940 1.400 1256.780 1279.600 ;
    RECT 1257.060 1.400 1257.900 1279.600 ;
    RECT 1258.180 1.400 1259.020 1279.600 ;
    RECT 1259.300 1.400 1260.140 1279.600 ;
    RECT 1260.420 1.400 1261.260 1279.600 ;
    RECT 1261.540 1.400 1262.380 1279.600 ;
    RECT 1262.660 1.400 1263.500 1279.600 ;
    RECT 1263.780 1.400 1264.620 1279.600 ;
    RECT 1264.900 1.400 1265.740 1279.600 ;
    RECT 1266.020 1.400 1266.860 1279.600 ;
    RECT 1267.140 1.400 1267.980 1279.600 ;
    RECT 1268.260 1.400 1269.100 1279.600 ;
    RECT 1269.380 1.400 1270.220 1279.600 ;
    RECT 1270.500 1.400 1271.340 1279.600 ;
    RECT 1271.620 1.400 1272.460 1279.600 ;
    RECT 1272.740 1.400 1273.580 1279.600 ;
    RECT 1273.860 1.400 1274.700 1279.600 ;
    RECT 1274.980 1.400 1275.820 1279.600 ;
    RECT 1276.100 1.400 1276.940 1279.600 ;
    RECT 1277.220 1.400 1278.060 1279.600 ;
    RECT 1278.340 1.400 1279.180 1279.600 ;
    RECT 1279.460 1.400 1280.300 1279.600 ;
    RECT 1280.580 1.400 1281.420 1279.600 ;
    RECT 1281.700 1.400 1282.540 1279.600 ;
    RECT 1282.820 1.400 1283.660 1279.600 ;
    RECT 1283.940 1.400 1284.780 1279.600 ;
    RECT 1285.060 1.400 1285.900 1279.600 ;
    RECT 1286.180 1.400 1287.020 1279.600 ;
    RECT 1287.300 1.400 1288.140 1279.600 ;
    RECT 1288.420 1.400 1289.260 1279.600 ;
    RECT 1289.540 1.400 1290.380 1279.600 ;
    RECT 1290.660 1.400 1291.500 1279.600 ;
    RECT 1291.780 1.400 1292.620 1279.600 ;
    RECT 1292.900 1.400 1293.740 1279.600 ;
    RECT 1294.020 1.400 1294.860 1279.600 ;
    RECT 1295.140 1.400 1295.980 1279.600 ;
    RECT 1296.260 1.400 1297.100 1279.600 ;
    RECT 1297.380 1.400 1298.220 1279.600 ;
    RECT 1298.500 1.400 1299.340 1279.600 ;
    RECT 1299.620 1.400 1300.460 1279.600 ;
    RECT 1300.740 1.400 1301.580 1279.600 ;
    RECT 1301.860 1.400 1302.700 1279.600 ;
    RECT 1302.980 1.400 1303.820 1279.600 ;
    RECT 1304.100 1.400 1304.940 1279.600 ;
    RECT 1305.220 1.400 1306.060 1279.600 ;
    RECT 1306.340 1.400 1307.180 1279.600 ;
    RECT 1307.460 1.400 1308.300 1279.600 ;
    RECT 1308.580 1.400 1309.420 1279.600 ;
    RECT 1309.700 1.400 1310.540 1279.600 ;
    RECT 1310.820 1.400 1311.660 1279.600 ;
    RECT 1311.940 1.400 1312.780 1279.600 ;
    RECT 1313.060 1.400 1313.900 1279.600 ;
    RECT 1314.180 1.400 1315.020 1279.600 ;
    RECT 1315.300 1.400 1316.140 1279.600 ;
    RECT 1316.420 1.400 1317.260 1279.600 ;
    RECT 1317.540 1.400 1318.380 1279.600 ;
    RECT 1318.660 1.400 1319.500 1279.600 ;
    RECT 1319.780 1.400 1320.620 1279.600 ;
    RECT 1320.900 1.400 1321.740 1279.600 ;
    RECT 1322.020 1.400 1322.860 1279.600 ;
    RECT 1323.140 1.400 1323.980 1279.600 ;
    RECT 1324.260 1.400 1325.100 1279.600 ;
    RECT 1325.380 1.400 1326.220 1279.600 ;
    RECT 1326.500 1.400 1327.340 1279.600 ;
    RECT 1327.620 1.400 1328.460 1279.600 ;
    RECT 1328.740 1.400 1329.580 1279.600 ;
    RECT 1329.860 1.400 1330.700 1279.600 ;
    RECT 1330.980 1.400 1331.820 1279.600 ;
    RECT 1332.100 1.400 1332.940 1279.600 ;
    RECT 1333.220 1.400 1334.060 1279.600 ;
    RECT 1334.340 1.400 1335.180 1279.600 ;
    RECT 1335.460 1.400 1336.300 1279.600 ;
    RECT 1336.580 1.400 1337.420 1279.600 ;
    RECT 1337.700 1.400 1338.540 1279.600 ;
    RECT 1338.820 1.400 1339.660 1279.600 ;
    RECT 1339.940 1.400 1340.780 1279.600 ;
    RECT 1341.060 1.400 1341.900 1279.600 ;
    RECT 1342.180 1.400 1343.020 1279.600 ;
    RECT 1343.300 1.400 1344.140 1279.600 ;
    RECT 1344.420 1.400 1345.260 1279.600 ;
    RECT 1345.540 1.400 1346.380 1279.600 ;
    RECT 1346.660 1.400 1347.500 1279.600 ;
    RECT 1347.780 1.400 1348.620 1279.600 ;
    RECT 1348.900 1.400 1349.740 1279.600 ;
    RECT 1350.020 1.400 1350.860 1279.600 ;
    RECT 1351.140 1.400 1351.980 1279.600 ;
    RECT 1352.260 1.400 1353.100 1279.600 ;
    RECT 1353.380 1.400 1354.220 1279.600 ;
    RECT 1354.500 1.400 1355.340 1279.600 ;
    RECT 1355.620 1.400 1356.460 1279.600 ;
    RECT 1356.740 1.400 1357.580 1279.600 ;
    RECT 1357.860 1.400 1358.700 1279.600 ;
    RECT 1358.980 1.400 1359.820 1279.600 ;
    RECT 1360.100 1.400 1360.940 1279.600 ;
    RECT 1361.220 1.400 1362.060 1279.600 ;
    RECT 1362.340 1.400 1363.180 1279.600 ;
    RECT 1363.460 1.400 1364.300 1279.600 ;
    RECT 1364.580 1.400 1365.420 1279.600 ;
    RECT 1365.700 1.400 1366.540 1279.600 ;
    RECT 1366.820 1.400 1367.660 1279.600 ;
    RECT 1367.940 1.400 1368.780 1279.600 ;
    RECT 1369.060 1.400 1369.900 1279.600 ;
    RECT 1370.180 1.400 1371.020 1279.600 ;
    RECT 1371.300 1.400 1372.140 1279.600 ;
    RECT 1372.420 1.400 1373.260 1279.600 ;
    RECT 1373.540 1.400 1374.380 1279.600 ;
    RECT 1374.660 1.400 1375.500 1279.600 ;
    RECT 1375.780 1.400 1376.620 1279.600 ;
    RECT 1376.900 1.400 1377.740 1279.600 ;
    RECT 1378.020 1.400 1378.860 1279.600 ;
    RECT 1379.140 1.400 1379.980 1279.600 ;
    RECT 1380.260 1.400 1381.100 1279.600 ;
    RECT 1381.380 1.400 1382.220 1279.600 ;
    RECT 1382.500 1.400 1383.340 1279.600 ;
    RECT 1383.620 1.400 1384.460 1279.600 ;
    RECT 1384.740 1.400 1385.580 1279.600 ;
    RECT 1385.860 1.400 1386.700 1279.600 ;
    RECT 1386.980 1.400 1387.820 1279.600 ;
    RECT 1388.100 1.400 1388.940 1279.600 ;
    RECT 1389.220 1.400 1390.060 1279.600 ;
    RECT 1390.340 1.400 1391.180 1279.600 ;
    RECT 1391.460 1.400 1392.300 1279.600 ;
    RECT 1392.580 1.400 1393.420 1279.600 ;
    RECT 1393.700 1.400 1394.540 1279.600 ;
    RECT 1394.820 1.400 1395.660 1279.600 ;
    RECT 1395.940 1.400 1396.780 1279.600 ;
    RECT 1397.060 1.400 1397.900 1279.600 ;
    RECT 1398.180 1.400 1399.020 1279.600 ;
    RECT 1399.300 1.400 1400.140 1279.600 ;
    RECT 1400.420 1.400 1401.260 1279.600 ;
    RECT 1401.540 1.400 1402.380 1279.600 ;
    RECT 1402.660 1.400 1403.500 1279.600 ;
    RECT 1403.780 1.400 1404.620 1279.600 ;
    RECT 1404.900 1.400 1405.740 1279.600 ;
    RECT 1406.020 1.400 1406.860 1279.600 ;
    RECT 1407.140 1.400 1407.980 1279.600 ;
    RECT 1408.260 1.400 1409.100 1279.600 ;
    RECT 1409.380 1.400 1410.220 1279.600 ;
    RECT 1410.500 1.400 1411.340 1279.600 ;
    RECT 1411.620 1.400 1412.460 1279.600 ;
    RECT 1412.740 1.400 1413.580 1279.600 ;
    RECT 1413.860 1.400 1414.700 1279.600 ;
    RECT 1414.980 1.400 1415.820 1279.600 ;
    RECT 1416.100 1.400 1416.940 1279.600 ;
    RECT 1417.220 1.400 1418.060 1279.600 ;
    RECT 1418.340 1.400 1419.180 1279.600 ;
    RECT 1419.460 1.400 1420.300 1279.600 ;
    RECT 1420.580 1.400 1421.420 1279.600 ;
    RECT 1421.700 1.400 1422.540 1279.600 ;
    RECT 1422.820 1.400 1423.660 1279.600 ;
    RECT 1423.940 1.400 1424.780 1279.600 ;
    RECT 1425.060 1.400 1425.900 1279.600 ;
    RECT 1426.180 1.400 1427.020 1279.600 ;
    RECT 1427.300 1.400 1428.140 1279.600 ;
    RECT 1428.420 1.400 1429.260 1279.600 ;
    RECT 1429.540 1.400 1430.380 1279.600 ;
    RECT 1430.660 1.400 1431.500 1279.600 ;
    RECT 1431.780 1.400 1432.620 1279.600 ;
    RECT 1432.900 1.400 1433.740 1279.600 ;
    RECT 1434.020 1.400 1434.860 1279.600 ;
    RECT 1435.140 1.400 1435.980 1279.600 ;
    RECT 1436.260 1.400 1437.100 1279.600 ;
    RECT 1437.380 1.400 1438.220 1279.600 ;
    RECT 1438.500 1.400 1439.340 1279.600 ;
    RECT 1439.620 1.400 1440.460 1279.600 ;
    RECT 1440.740 1.400 1441.580 1279.600 ;
    RECT 1441.860 1.400 1442.700 1279.600 ;
    RECT 1442.980 1.400 1443.820 1279.600 ;
    RECT 1444.100 1.400 1444.940 1279.600 ;
    RECT 1445.220 1.400 1446.060 1279.600 ;
    RECT 1446.340 1.400 1447.180 1279.600 ;
    RECT 1447.460 1.400 1448.300 1279.600 ;
    RECT 1448.580 1.400 1449.420 1279.600 ;
    RECT 1449.700 1.400 1450.540 1279.600 ;
    RECT 1450.820 1.400 1451.660 1279.600 ;
    RECT 1451.940 1.400 1452.780 1279.600 ;
    RECT 1453.060 1.400 1453.900 1279.600 ;
    RECT 1454.180 1.400 1455.020 1279.600 ;
    RECT 1455.300 1.400 1456.140 1279.600 ;
    RECT 1456.420 1.400 1457.260 1279.600 ;
    RECT 1457.540 1.400 1458.380 1279.600 ;
    RECT 1458.660 1.400 1459.500 1279.600 ;
    RECT 1459.780 1.400 1460.620 1279.600 ;
    RECT 1460.900 1.400 1461.740 1279.600 ;
    RECT 1462.020 1.400 1462.860 1279.600 ;
    RECT 1463.140 1.400 1463.980 1279.600 ;
    RECT 1464.260 1.400 1465.100 1279.600 ;
    RECT 1465.380 1.400 1466.220 1279.600 ;
    RECT 1466.500 1.400 1467.340 1279.600 ;
    RECT 1467.620 1.400 1468.460 1279.600 ;
    RECT 1468.740 1.400 1469.580 1279.600 ;
    RECT 1469.860 1.400 1470.700 1279.600 ;
    RECT 1470.980 1.400 1471.820 1279.600 ;
    RECT 1472.100 1.400 1472.940 1279.600 ;
    RECT 1473.220 1.400 1474.060 1279.600 ;
    RECT 1474.340 1.400 1475.180 1279.600 ;
    RECT 1475.460 1.400 1476.300 1279.600 ;
    RECT 1476.580 1.400 1477.420 1279.600 ;
    RECT 1477.700 1.400 1478.540 1279.600 ;
    RECT 1478.820 1.400 1479.660 1279.600 ;
    RECT 1479.940 1.400 1480.780 1279.600 ;
    RECT 1481.060 1.400 1481.900 1279.600 ;
    RECT 1482.180 1.400 1483.020 1279.600 ;
    RECT 1483.300 1.400 1484.140 1279.600 ;
    RECT 1484.420 1.400 1485.260 1279.600 ;
    RECT 1485.540 1.400 1486.380 1279.600 ;
    RECT 1486.660 1.400 1487.500 1279.600 ;
    RECT 1487.780 1.400 1488.620 1279.600 ;
    RECT 1488.900 1.400 1489.740 1279.600 ;
    RECT 1490.020 1.400 1490.860 1279.600 ;
    RECT 1491.140 1.400 1491.980 1279.600 ;
    RECT 1492.260 1.400 1493.100 1279.600 ;
    RECT 1493.380 1.400 1494.220 1279.600 ;
    RECT 1494.500 1.400 1495.340 1279.600 ;
    RECT 1495.620 1.400 1496.460 1279.600 ;
    RECT 1496.740 1.400 1497.580 1279.600 ;
    RECT 1497.860 1.400 1498.700 1279.600 ;
    RECT 1498.980 1.400 1499.820 1279.600 ;
    RECT 1500.100 1.400 1500.940 1279.600 ;
    RECT 1501.220 1.400 1502.060 1279.600 ;
    RECT 1502.340 1.400 1503.180 1279.600 ;
    RECT 1503.460 1.400 1504.300 1279.600 ;
    RECT 1504.580 1.400 1505.420 1279.600 ;
    RECT 1505.700 1.400 1506.540 1279.600 ;
    RECT 1506.820 1.400 1507.660 1279.600 ;
    RECT 1507.940 1.400 1508.780 1279.600 ;
    RECT 1509.060 1.400 1509.900 1279.600 ;
    RECT 1510.180 1.400 1511.020 1279.600 ;
    RECT 1511.300 1.400 1512.140 1279.600 ;
    RECT 1512.420 1.400 1513.260 1279.600 ;
    RECT 1513.540 1.400 1514.380 1279.600 ;
    RECT 1514.660 1.400 1515.500 1279.600 ;
    RECT 1515.780 1.400 1516.620 1279.600 ;
    RECT 1516.900 1.400 1517.740 1279.600 ;
    RECT 1518.020 1.400 1518.860 1279.600 ;
    RECT 1519.140 1.400 1519.980 1279.600 ;
    RECT 1520.260 1.400 1521.100 1279.600 ;
    RECT 1521.380 1.400 1522.220 1279.600 ;
    RECT 1522.500 1.400 1523.340 1279.600 ;
    RECT 1523.620 1.400 1524.460 1279.600 ;
    RECT 1524.740 1.400 1525.580 1279.600 ;
    RECT 1525.860 1.400 1526.700 1279.600 ;
    RECT 1526.980 1.400 1527.820 1279.600 ;
    RECT 1528.100 1.400 1528.940 1279.600 ;
    RECT 1529.220 1.400 1530.060 1279.600 ;
    RECT 1530.340 1.400 1531.180 1279.600 ;
    RECT 1531.460 1.400 1532.300 1279.600 ;
    RECT 1532.580 1.400 1533.420 1279.600 ;
    RECT 1533.700 1.400 1534.540 1279.600 ;
    RECT 1534.820 1.400 1535.660 1279.600 ;
    RECT 1535.940 1.400 1536.780 1279.600 ;
    RECT 1537.060 1.400 1537.900 1279.600 ;
    RECT 1538.180 1.400 1539.020 1279.600 ;
    RECT 1539.300 1.400 1540.140 1279.600 ;
    RECT 1540.420 1.400 1541.260 1279.600 ;
    RECT 1541.540 1.400 1542.380 1279.600 ;
    RECT 1542.660 1.400 1543.500 1279.600 ;
    RECT 1543.780 1.400 1544.620 1279.600 ;
    RECT 1544.900 1.400 1545.740 1279.600 ;
    RECT 1546.020 1.400 1546.860 1279.600 ;
    RECT 1547.140 1.400 1547.980 1279.600 ;
    RECT 1548.260 1.400 1549.100 1279.600 ;
    RECT 1549.380 1.400 1550.220 1279.600 ;
    RECT 1550.500 1.400 1551.340 1279.600 ;
    RECT 1551.620 1.400 1552.460 1279.600 ;
    RECT 1552.740 1.400 1553.580 1279.600 ;
    RECT 1553.860 1.400 1554.700 1279.600 ;
    RECT 1554.980 1.400 1555.820 1279.600 ;
    RECT 1556.100 1.400 1556.940 1279.600 ;
    RECT 1557.220 1.400 1558.060 1279.600 ;
    RECT 1558.340 1.400 1559.180 1279.600 ;
    RECT 1559.460 1.400 1560.300 1279.600 ;
    RECT 1560.580 1.400 1561.420 1279.600 ;
    RECT 1561.700 1.400 1562.540 1279.600 ;
    RECT 1562.820 1.400 1563.660 1279.600 ;
    RECT 1563.940 1.400 1564.780 1279.600 ;
    RECT 1565.060 1.400 1565.900 1279.600 ;
    RECT 1566.180 1.400 1567.020 1279.600 ;
    RECT 1567.300 1.400 1568.140 1279.600 ;
    RECT 1568.420 1.400 1569.260 1279.600 ;
    RECT 1569.540 1.400 1570.380 1279.600 ;
    RECT 1570.660 1.400 1571.500 1279.600 ;
    RECT 1571.780 1.400 1572.620 1279.600 ;
    RECT 1572.900 1.400 1573.740 1279.600 ;
    RECT 1574.020 1.400 1574.860 1279.600 ;
    RECT 1575.140 1.400 1575.980 1279.600 ;
    RECT 1576.260 1.400 1577.100 1279.600 ;
    RECT 1577.380 1.400 1578.220 1279.600 ;
    RECT 1578.500 1.400 1579.340 1279.600 ;
    RECT 1579.620 1.400 1580.460 1279.600 ;
    RECT 1580.740 1.400 1581.580 1279.600 ;
    RECT 1581.860 1.400 1582.700 1279.600 ;
    RECT 1582.980 1.400 1583.820 1279.600 ;
    RECT 1584.100 1.400 1584.940 1279.600 ;
    RECT 1585.220 1.400 1586.060 1279.600 ;
    RECT 1586.340 1.400 1587.180 1279.600 ;
    RECT 1587.460 1.400 1588.300 1279.600 ;
    RECT 1588.580 1.400 1589.420 1279.600 ;
    RECT 1589.700 1.400 1590.540 1279.600 ;
    RECT 1590.820 1.400 1591.660 1279.600 ;
    RECT 1591.940 1.400 1592.780 1279.600 ;
    RECT 1593.060 1.400 1593.900 1279.600 ;
    RECT 1594.180 1.400 1595.020 1279.600 ;
    RECT 1595.300 1.400 1596.140 1279.600 ;
    RECT 1596.420 1.400 1597.260 1279.600 ;
    RECT 1597.540 1.400 1598.380 1279.600 ;
    RECT 1598.660 1.400 1599.500 1279.600 ;
    RECT 1599.780 1.400 1600.620 1279.600 ;
    RECT 1600.900 1.400 1601.740 1279.600 ;
    RECT 1602.020 1.400 1602.860 1279.600 ;
    RECT 1603.140 1.400 1603.980 1279.600 ;
    RECT 1604.260 1.400 1605.100 1279.600 ;
    RECT 1605.380 1.400 1606.220 1279.600 ;
    RECT 1606.500 1.400 1607.340 1279.600 ;
    RECT 1607.620 1.400 1608.460 1279.600 ;
    RECT 1608.740 1.400 1609.580 1279.600 ;
    RECT 1609.860 1.400 1610.700 1279.600 ;
    RECT 1610.980 1.400 1611.820 1279.600 ;
    RECT 1612.100 1.400 1612.940 1279.600 ;
    RECT 1613.220 1.400 1614.060 1279.600 ;
    RECT 1614.340 1.400 1615.180 1279.600 ;
    RECT 1615.460 1.400 1616.300 1279.600 ;
    RECT 1616.580 1.400 1617.420 1279.600 ;
    RECT 1617.700 1.400 1618.540 1279.600 ;
    RECT 1618.820 1.400 1619.660 1279.600 ;
    RECT 1619.940 1.400 1620.780 1279.600 ;
    RECT 1621.060 1.400 1621.900 1279.600 ;
    RECT 1622.180 1.400 1623.020 1279.600 ;
    RECT 1623.300 1.400 1624.140 1279.600 ;
    RECT 1624.420 1.400 1625.260 1279.600 ;
    RECT 1625.540 1.400 1626.380 1279.600 ;
    RECT 1626.660 1.400 1627.500 1279.600 ;
    RECT 1627.780 1.400 1628.620 1279.600 ;
    RECT 1628.900 1.400 1629.740 1279.600 ;
    RECT 1630.020 1.400 1630.860 1279.600 ;
    RECT 1631.140 1.400 1631.980 1279.600 ;
    RECT 1632.260 1.400 1633.100 1279.600 ;
    RECT 1633.380 1.400 1634.220 1279.600 ;
    RECT 1634.500 1.400 1635.340 1279.600 ;
    RECT 1635.620 1.400 1636.460 1279.600 ;
    RECT 1636.740 1.400 1637.580 1279.600 ;
    RECT 1637.860 1.400 1638.700 1279.600 ;
    RECT 1638.980 1.400 1639.820 1279.600 ;
    RECT 1640.100 1.400 1640.940 1279.600 ;
    RECT 1641.220 1.400 1642.060 1279.600 ;
    RECT 1642.340 1.400 1643.180 1279.600 ;
    RECT 1643.460 1.400 1644.300 1279.600 ;
    RECT 1644.580 1.400 1645.420 1279.600 ;
    RECT 1645.700 1.400 1646.540 1279.600 ;
    RECT 1646.820 1.400 1647.660 1279.600 ;
    RECT 1647.940 1.400 1648.780 1279.600 ;
    RECT 1649.060 1.400 1649.900 1279.600 ;
    RECT 1650.180 1.400 1651.020 1279.600 ;
    RECT 1651.300 1.400 1652.140 1279.600 ;
    RECT 1652.420 1.400 1653.260 1279.600 ;
    RECT 1653.540 1.400 1654.380 1279.600 ;
    RECT 1654.660 1.400 1655.500 1279.600 ;
    RECT 1655.780 1.400 1656.620 1279.600 ;
    RECT 1656.900 1.400 1657.740 1279.600 ;
    RECT 1658.020 1.400 1658.860 1279.600 ;
    RECT 1659.140 1.400 1659.980 1279.600 ;
    RECT 1660.260 1.400 1661.100 1279.600 ;
    RECT 1661.380 1.400 1662.220 1279.600 ;
    RECT 1662.500 1.400 1663.340 1279.600 ;
    RECT 1663.620 1.400 1664.460 1279.600 ;
    RECT 1664.740 1.400 1665.580 1279.600 ;
    RECT 1665.860 1.400 1666.700 1279.600 ;
    RECT 1666.980 1.400 1667.820 1279.600 ;
    RECT 1668.100 1.400 1668.940 1279.600 ;
    RECT 1669.220 1.400 1670.060 1279.600 ;
    RECT 1670.340 1.400 1671.180 1279.600 ;
    RECT 1671.460 1.400 1672.300 1279.600 ;
    RECT 1672.580 1.400 1673.420 1279.600 ;
    RECT 1673.700 1.400 1674.540 1279.600 ;
    RECT 1674.820 1.400 1675.660 1279.600 ;
    RECT 1675.940 1.400 1676.780 1279.600 ;
    RECT 1677.060 1.400 1677.900 1279.600 ;
    RECT 1678.180 1.400 1679.020 1279.600 ;
    RECT 1679.300 1.400 1680.140 1279.600 ;
    RECT 1680.420 1.400 1681.260 1279.600 ;
    RECT 1681.540 1.400 1682.380 1279.600 ;
    RECT 1682.660 1.400 1683.500 1279.600 ;
    RECT 1683.780 1.400 1684.620 1279.600 ;
    RECT 1684.900 1.400 1685.740 1279.600 ;
    RECT 1686.020 1.400 1686.860 1279.600 ;
    RECT 1687.140 1.400 1687.980 1279.600 ;
    RECT 1688.260 1.400 1689.100 1279.600 ;
    RECT 1689.380 1.400 1690.220 1279.600 ;
    RECT 1690.500 1.400 1691.340 1279.600 ;
    RECT 1691.620 1.400 1692.460 1279.600 ;
    RECT 1692.740 1.400 1693.580 1279.600 ;
    RECT 1693.860 1.400 1694.700 1279.600 ;
    RECT 1694.980 1.400 1695.820 1279.600 ;
    RECT 1696.100 1.400 1696.940 1279.600 ;
    RECT 1697.220 1.400 1698.060 1279.600 ;
    RECT 1698.340 1.400 1699.180 1279.600 ;
    RECT 1699.460 1.400 1700.300 1279.600 ;
    RECT 1700.580 1.400 1701.420 1279.600 ;
    RECT 1701.700 1.400 1702.540 1279.600 ;
    RECT 1702.820 1.400 1703.660 1279.600 ;
    RECT 1703.940 1.400 1704.780 1279.600 ;
    RECT 1705.060 1.400 1705.900 1279.600 ;
    RECT 1706.180 1.400 1707.020 1279.600 ;
    RECT 1707.300 1.400 1708.140 1279.600 ;
    RECT 1708.420 1.400 1709.260 1279.600 ;
    RECT 1709.540 1.400 1710.380 1279.600 ;
    RECT 1710.660 1.400 1711.500 1279.600 ;
    RECT 1711.780 1.400 1712.620 1279.600 ;
    RECT 1712.900 1.400 1713.740 1279.600 ;
    RECT 1714.020 1.400 1714.860 1279.600 ;
    RECT 1715.140 1.400 1715.980 1279.600 ;
    RECT 1716.260 1.400 1717.100 1279.600 ;
    RECT 1717.380 1.400 1718.220 1279.600 ;
    RECT 1718.500 1.400 1719.340 1279.600 ;
    RECT 1719.620 1.400 1720.460 1279.600 ;
    RECT 1720.740 1.400 1721.580 1279.600 ;
    RECT 1721.860 1.400 1722.700 1279.600 ;
    RECT 1722.980 1.400 1723.820 1279.600 ;
    RECT 1724.100 1.400 1724.940 1279.600 ;
    RECT 1725.220 1.400 1726.060 1279.600 ;
    RECT 1726.340 1.400 1727.180 1279.600 ;
    RECT 1727.460 1.400 1728.300 1279.600 ;
    RECT 1728.580 1.400 1729.420 1279.600 ;
    RECT 1729.700 1.400 1730.540 1279.600 ;
    RECT 1730.820 1.400 1731.660 1279.600 ;
    RECT 1731.940 1.400 1732.780 1279.600 ;
    RECT 1733.060 1.400 1733.900 1279.600 ;
    RECT 1734.180 1.400 1735.020 1279.600 ;
    RECT 1735.300 1.400 1736.140 1279.600 ;
    RECT 1736.420 1.400 1737.260 1279.600 ;
    RECT 1737.540 1.400 1738.380 1279.600 ;
    RECT 1738.660 1.400 1739.500 1279.600 ;
    RECT 1739.780 1.400 1740.620 1279.600 ;
    RECT 1740.900 1.400 1741.740 1279.600 ;
    RECT 1742.020 1.400 1742.860 1279.600 ;
    RECT 1743.140 1.400 1743.980 1279.600 ;
    RECT 1744.260 1.400 1745.100 1279.600 ;
    RECT 1745.380 1.400 1746.220 1279.600 ;
    RECT 1746.500 1.400 1747.340 1279.600 ;
    RECT 1747.620 1.400 1748.460 1279.600 ;
    RECT 1748.740 1.400 1749.580 1279.600 ;
    RECT 1749.860 1.400 1750.700 1279.600 ;
    RECT 1750.980 1.400 1751.820 1279.600 ;
    RECT 1752.100 1.400 1752.940 1279.600 ;
    RECT 1753.220 1.400 1754.060 1279.600 ;
    RECT 1754.340 1.400 1755.180 1279.600 ;
    RECT 1755.460 1.400 1756.300 1279.600 ;
    RECT 1756.580 1.400 1757.420 1279.600 ;
    RECT 1757.700 1.400 1758.540 1279.600 ;
    RECT 1758.820 1.400 1759.660 1279.600 ;
    RECT 1759.940 1.400 1760.780 1279.600 ;
    RECT 1761.060 1.400 1761.900 1279.600 ;
    RECT 1762.180 1.400 1763.020 1279.600 ;
    RECT 1763.300 1.400 1764.140 1279.600 ;
    RECT 1764.420 1.400 1765.260 1279.600 ;
    RECT 1765.540 1.400 1766.380 1279.600 ;
    RECT 1766.660 1.400 1767.500 1279.600 ;
    RECT 1767.780 1.400 1768.620 1279.600 ;
    RECT 1768.900 1.400 1769.740 1279.600 ;
    RECT 1770.020 1.400 1770.860 1279.600 ;
    RECT 1771.140 1.400 1771.980 1279.600 ;
    RECT 1772.260 1.400 1773.100 1279.600 ;
    RECT 1773.380 1.400 1774.220 1279.600 ;
    RECT 1774.500 1.400 1775.340 1279.600 ;
    RECT 1775.620 1.400 1776.460 1279.600 ;
    RECT 1776.740 1.400 1777.580 1279.600 ;
    RECT 1777.860 1.400 1778.700 1279.600 ;
    RECT 1778.980 1.400 1779.820 1279.600 ;
    RECT 1780.100 1.400 1780.940 1279.600 ;
    RECT 1781.220 1.400 1782.060 1279.600 ;
    RECT 1782.340 1.400 1783.180 1279.600 ;
    RECT 1783.460 1.400 1784.300 1279.600 ;
    RECT 1784.580 1.400 1785.420 1279.600 ;
    RECT 1785.700 1.400 1786.540 1279.600 ;
    RECT 1786.820 1.400 1787.660 1279.600 ;
    RECT 1787.940 1.400 1788.780 1279.600 ;
    RECT 1789.060 1.400 1789.900 1279.600 ;
    RECT 1790.180 1.400 1791.020 1279.600 ;
    RECT 1791.300 1.400 1792.140 1279.600 ;
    RECT 1792.420 1.400 1793.260 1279.600 ;
    RECT 1793.540 1.400 1794.380 1279.600 ;
    RECT 1794.660 1.400 1795.500 1279.600 ;
    RECT 1795.780 1.400 1796.620 1279.600 ;
    RECT 1796.900 1.400 1797.740 1279.600 ;
    RECT 1798.020 1.400 1798.860 1279.600 ;
    RECT 1799.140 1.400 1799.980 1279.600 ;
    RECT 1800.260 1.400 1801.100 1279.600 ;
    RECT 1801.380 1.400 1802.220 1279.600 ;
    RECT 1802.500 1.400 1803.340 1279.600 ;
    RECT 1803.620 1.400 1804.460 1279.600 ;
    RECT 1804.740 1.400 1805.580 1279.600 ;
    RECT 1805.860 1.400 1806.700 1279.600 ;
    RECT 1806.980 1.400 1807.820 1279.600 ;
    RECT 1808.100 1.400 1808.940 1279.600 ;
    RECT 1809.220 1.400 1810.060 1279.600 ;
    RECT 1810.340 1.400 1811.180 1279.600 ;
    RECT 1811.460 1.400 1812.300 1279.600 ;
    RECT 1812.580 1.400 1813.420 1279.600 ;
    RECT 1813.700 1.400 1814.540 1279.600 ;
    RECT 1814.820 1.400 1815.660 1279.600 ;
    RECT 1815.940 1.400 1816.780 1279.600 ;
    RECT 1817.060 1.400 1817.900 1279.600 ;
    RECT 1818.180 1.400 1819.020 1279.600 ;
    RECT 1819.300 1.400 1820.140 1279.600 ;
    RECT 1820.420 1.400 1821.260 1279.600 ;
    RECT 1821.540 1.400 1822.380 1279.600 ;
    RECT 1822.660 1.400 1823.500 1279.600 ;
    RECT 1823.780 1.400 1824.620 1279.600 ;
    RECT 1824.900 1.400 1825.740 1279.600 ;
    RECT 1826.020 1.400 1826.860 1279.600 ;
    RECT 1827.140 1.400 1827.980 1279.600 ;
    RECT 1828.260 1.400 1829.100 1279.600 ;
    RECT 1829.380 1.400 1830.220 1279.600 ;
    RECT 1830.500 1.400 1831.340 1279.600 ;
    RECT 1831.620 1.400 1832.460 1279.600 ;
    RECT 1832.740 1.400 1833.580 1279.600 ;
    RECT 1833.860 1.400 1834.700 1279.600 ;
    RECT 1834.980 1.400 1835.820 1279.600 ;
    RECT 1836.100 1.400 1836.940 1279.600 ;
    RECT 1837.220 1.400 1838.060 1279.600 ;
    RECT 1838.340 1.400 1839.180 1279.600 ;
    RECT 1839.460 1.400 1840.300 1279.600 ;
    RECT 1840.580 1.400 1841.420 1279.600 ;
    RECT 1841.700 1.400 1842.540 1279.600 ;
    RECT 1842.820 1.400 1843.660 1279.600 ;
    RECT 1843.940 1.400 1844.780 1279.600 ;
    RECT 1845.060 1.400 1845.900 1279.600 ;
    RECT 1846.180 1.400 1847.020 1279.600 ;
    RECT 1847.300 1.400 1848.140 1279.600 ;
    RECT 1848.420 1.400 1849.260 1279.600 ;
    RECT 1849.540 1.400 1850.380 1279.600 ;
    RECT 1850.660 1.400 1851.500 1279.600 ;
    RECT 1851.780 1.400 1852.620 1279.600 ;
    RECT 1852.900 1.400 1853.740 1279.600 ;
    RECT 1854.020 1.400 1854.860 1279.600 ;
    RECT 1855.140 1.400 1855.980 1279.600 ;
    RECT 1856.260 1.400 1857.100 1279.600 ;
    RECT 1857.380 1.400 1858.220 1279.600 ;
    RECT 1858.500 1.400 1859.340 1279.600 ;
    RECT 1859.620 1.400 1860.460 1279.600 ;
    RECT 1860.740 1.400 1861.580 1279.600 ;
    RECT 1861.860 1.400 1862.700 1279.600 ;
    RECT 1862.980 1.400 1863.820 1279.600 ;
    RECT 1864.100 1.400 1864.940 1279.600 ;
    RECT 1865.220 1.400 1866.060 1279.600 ;
    RECT 1866.340 1.400 1867.180 1279.600 ;
    RECT 1867.460 1.400 1868.300 1279.600 ;
    RECT 1868.580 1.400 1869.420 1279.600 ;
    RECT 1869.700 1.400 1870.540 1279.600 ;
    RECT 1870.820 1.400 1871.660 1279.600 ;
    RECT 1871.940 1.400 1872.780 1279.600 ;
    RECT 1873.060 1.400 1873.900 1279.600 ;
    RECT 1874.180 1.400 1875.020 1279.600 ;
    RECT 1875.300 1.400 1876.140 1279.600 ;
    RECT 1876.420 1.400 1877.260 1279.600 ;
    RECT 1877.540 1.400 1878.380 1279.600 ;
    RECT 1878.660 1.400 1879.500 1279.600 ;
    RECT 1879.780 1.400 1880.620 1279.600 ;
    RECT 1880.900 1.400 1881.740 1279.600 ;
    RECT 1882.020 1.400 1882.860 1279.600 ;
    RECT 1883.140 1.400 1883.980 1279.600 ;
    RECT 1884.260 1.400 1885.100 1279.600 ;
    RECT 1885.380 1.400 1886.220 1279.600 ;
    RECT 1886.500 1.400 1887.340 1279.600 ;
    RECT 1887.620 1.400 1888.460 1279.600 ;
    RECT 1888.740 1.400 1889.580 1279.600 ;
    RECT 1889.860 1.400 1890.700 1279.600 ;
    RECT 1890.980 1.400 1891.820 1279.600 ;
    RECT 1892.100 1.400 1892.940 1279.600 ;
    RECT 1893.220 1.400 1894.060 1279.600 ;
    RECT 1894.340 1.400 1895.180 1279.600 ;
    RECT 1895.460 1.400 1896.300 1279.600 ;
    RECT 1896.580 1.400 1897.420 1279.600 ;
    RECT 1897.700 1.400 1898.540 1279.600 ;
    RECT 1898.820 1.400 1899.660 1279.600 ;
    RECT 1899.940 1.400 1900.780 1279.600 ;
    RECT 1901.060 1.400 1901.900 1279.600 ;
    RECT 1902.180 1.400 1903.020 1279.600 ;
    RECT 1903.300 1.400 1904.140 1279.600 ;
    RECT 1904.420 1.400 1905.260 1279.600 ;
    RECT 1905.540 1.400 1906.380 1279.600 ;
    RECT 1906.660 1.400 1907.500 1279.600 ;
    RECT 1907.780 1.400 1908.620 1279.600 ;
    RECT 1908.900 1.400 1909.740 1279.600 ;
    RECT 1910.020 1.400 1910.860 1279.600 ;
    RECT 1911.140 1.400 1911.980 1279.600 ;
    RECT 1912.260 1.400 1913.100 1279.600 ;
    RECT 1913.380 1.400 1914.220 1279.600 ;
    RECT 1914.500 1.400 1915.340 1279.600 ;
    RECT 1915.620 1.400 1916.460 1279.600 ;
    RECT 1916.740 1.400 1917.580 1279.600 ;
    RECT 1917.860 1.400 1918.700 1279.600 ;
    RECT 1918.980 1.400 1919.820 1279.600 ;
    RECT 1920.100 1.400 1920.940 1279.600 ;
    RECT 1921.220 1.400 1922.060 1279.600 ;
    RECT 1922.340 1.400 1923.180 1279.600 ;
    RECT 1923.460 1.400 1924.300 1279.600 ;
    RECT 1924.580 1.400 1925.420 1279.600 ;
    RECT 1925.700 1.400 1926.540 1279.600 ;
    RECT 1926.820 1.400 1927.660 1279.600 ;
    RECT 1927.940 1.400 1928.780 1279.600 ;
    RECT 1929.060 1.400 1929.900 1279.600 ;
    RECT 1930.180 1.400 1931.020 1279.600 ;
    RECT 1931.300 1.400 1932.140 1279.600 ;
    RECT 1932.420 1.400 1933.260 1279.600 ;
    RECT 1933.540 1.400 1934.380 1279.600 ;
    RECT 1934.660 1.400 1935.500 1279.600 ;
    RECT 1935.780 1.400 1936.620 1279.600 ;
    RECT 1936.900 1.400 1937.740 1279.600 ;
    RECT 1938.020 1.400 1938.860 1279.600 ;
    RECT 1939.140 1.400 1939.980 1279.600 ;
    RECT 1940.260 1.400 1941.100 1279.600 ;
    RECT 1941.380 1.400 1942.220 1279.600 ;
    RECT 1942.500 1.400 1943.340 1279.600 ;
    RECT 1943.620 1.400 1944.460 1279.600 ;
    RECT 1944.740 1.400 1945.580 1279.600 ;
    RECT 1945.860 1.400 1946.700 1279.600 ;
    RECT 1946.980 1.400 1947.820 1279.600 ;
    RECT 1948.100 1.400 1948.940 1279.600 ;
    RECT 1949.220 1.400 1950.060 1279.600 ;
    RECT 1950.340 1.400 1951.180 1279.600 ;
    RECT 1951.460 1.400 1952.300 1279.600 ;
    RECT 1952.580 1.400 1953.420 1279.600 ;
    RECT 1953.700 1.400 1954.540 1279.600 ;
    RECT 1954.820 1.400 1955.660 1279.600 ;
    RECT 1955.940 1.400 1956.780 1279.600 ;
    RECT 1957.060 1.400 1957.900 1279.600 ;
    RECT 1958.180 1.400 1959.020 1279.600 ;
    RECT 1959.300 1.400 1960.140 1279.600 ;
    RECT 1960.420 1.400 1961.260 1279.600 ;
    RECT 1961.540 1.400 1962.380 1279.600 ;
    RECT 1962.660 1.400 1963.500 1279.600 ;
    RECT 1963.780 1.400 1964.620 1279.600 ;
    RECT 1964.900 1.400 1965.740 1279.600 ;
    RECT 1966.020 1.400 1966.860 1279.600 ;
    RECT 1967.140 1.400 1967.980 1279.600 ;
    RECT 1968.260 1.400 1969.100 1279.600 ;
    RECT 1969.380 1.400 1970.220 1279.600 ;
    RECT 1970.500 1.400 1971.340 1279.600 ;
    RECT 1971.620 1.400 1972.460 1279.600 ;
    RECT 1972.740 1.400 1973.580 1279.600 ;
    RECT 1973.860 1.400 1974.700 1279.600 ;
    RECT 1974.980 1.400 1975.820 1279.600 ;
    RECT 1976.100 1.400 1976.940 1279.600 ;
    RECT 1977.220 1.400 1978.060 1279.600 ;
    RECT 1978.340 1.400 1979.180 1279.600 ;
    RECT 1979.460 1.400 1980.300 1279.600 ;
    RECT 1980.580 1.400 1981.420 1279.600 ;
    RECT 1981.700 1.400 1982.540 1279.600 ;
    RECT 1982.820 1.400 1983.660 1279.600 ;
    RECT 1983.940 1.400 1984.780 1279.600 ;
    RECT 1985.060 1.400 1985.900 1279.600 ;
    RECT 1986.180 1.400 1987.020 1279.600 ;
    RECT 1987.300 1.400 1988.140 1279.600 ;
    RECT 1988.420 1.400 1989.260 1279.600 ;
    RECT 1989.540 1.400 1990.380 1279.600 ;
    RECT 1990.660 1.400 1991.500 1279.600 ;
    RECT 1991.780 1.400 1992.620 1279.600 ;
    RECT 1992.900 1.400 1993.740 1279.600 ;
    RECT 1994.020 1.400 1994.860 1279.600 ;
    RECT 1995.140 1.400 1995.980 1279.600 ;
    RECT 1996.260 1.400 1997.100 1279.600 ;
    RECT 1997.380 1.400 1998.220 1279.600 ;
    RECT 1998.500 1.400 1999.340 1279.600 ;
    RECT 1999.620 1.400 2000.460 1279.600 ;
    RECT 2000.740 1.400 2001.580 1279.600 ;
    RECT 2001.860 1.400 2002.700 1279.600 ;
    RECT 2002.980 1.400 2003.820 1279.600 ;
    RECT 2004.100 1.400 2004.940 1279.600 ;
    RECT 2005.220 1.400 2006.060 1279.600 ;
    RECT 2006.340 1.400 2007.180 1279.600 ;
    RECT 2007.460 1.400 2008.300 1279.600 ;
    RECT 2008.580 1.400 2009.420 1279.600 ;
    RECT 2009.700 1.400 2010.540 1279.600 ;
    RECT 2010.820 1.400 2011.660 1279.600 ;
    RECT 2011.940 1.400 2012.780 1279.600 ;
    RECT 2013.060 1.400 2013.900 1279.600 ;
    RECT 2014.180 1.400 2015.020 1279.600 ;
    RECT 2015.300 1.400 2016.140 1279.600 ;
    RECT 2016.420 1.400 2017.260 1279.600 ;
    RECT 2017.540 1.400 2018.380 1279.600 ;
    RECT 2018.660 1.400 2019.500 1279.600 ;
    RECT 2019.780 1.400 2020.620 1279.600 ;
    RECT 2020.900 1.400 2021.740 1279.600 ;
    RECT 2022.020 1.400 2022.860 1279.600 ;
    RECT 2023.140 1.400 2023.980 1279.600 ;
    RECT 2024.260 1.400 2025.100 1279.600 ;
    RECT 2025.380 1.400 2026.220 1279.600 ;
    RECT 2026.500 1.400 2027.340 1279.600 ;
    RECT 2027.620 1.400 2028.460 1279.600 ;
    RECT 2028.740 1.400 2029.580 1279.600 ;
    RECT 2029.860 1.400 2030.700 1279.600 ;
    RECT 2030.980 1.400 2031.820 1279.600 ;
    RECT 2032.100 1.400 2032.940 1279.600 ;
    RECT 2033.220 1.400 2034.060 1279.600 ;
    RECT 2034.340 1.400 2035.180 1279.600 ;
    RECT 2035.460 1.400 2036.300 1279.600 ;
    RECT 2036.580 1.400 2037.420 1279.600 ;
    RECT 2037.700 1.400 2038.540 1279.600 ;
    RECT 2038.820 1.400 2039.660 1279.600 ;
    RECT 2039.940 1.400 2040.780 1279.600 ;
    RECT 2041.060 1.400 2041.900 1279.600 ;
    RECT 2042.180 1.400 2043.020 1279.600 ;
    RECT 2043.300 1.400 2044.140 1279.600 ;
    RECT 2044.420 1.400 2045.260 1279.600 ;
    RECT 2045.540 1.400 2046.380 1279.600 ;
    RECT 2046.660 1.400 2047.500 1279.600 ;
    RECT 2047.780 1.400 2048.620 1279.600 ;
    RECT 2048.900 1.400 2049.740 1279.600 ;
    RECT 2050.020 1.400 2050.860 1279.600 ;
    RECT 2051.140 1.400 2051.980 1279.600 ;
    RECT 2052.260 1.400 2053.100 1279.600 ;
    RECT 2053.380 1.400 2054.220 1279.600 ;
    RECT 2054.500 1.400 2055.340 1279.600 ;
    RECT 2055.620 1.400 2056.460 1279.600 ;
    RECT 2056.740 1.400 2057.580 1279.600 ;
    RECT 2057.860 1.400 2058.700 1279.600 ;
    RECT 2058.980 1.400 2059.820 1279.600 ;
    RECT 2060.100 1.400 2060.940 1279.600 ;
    RECT 2061.220 1.400 2062.060 1279.600 ;
    RECT 2062.340 1.400 2064.540 1279.600 ;
    LAYER OVERLAP ;
    RECT 0 0 2064.540 1281.000 ;
  END
END sram_512x4096_1rw

END LIBRARY
