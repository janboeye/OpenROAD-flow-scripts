VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_32x16384_1rw
  FOREIGN sram_32x16384_1rw 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1010.230 BY 616.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.805 0.070 91.875 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.125 0.070 97.195 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.765 0.070 107.835 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.405 0.070 118.475 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.725 0.070 123.795 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.045 0.070 129.115 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.365 0.070 134.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.685 0.070 139.755 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.645 0.070 155.715 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.965 0.070 161.035 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.285 0.070 166.355 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.225 0.070 169.295 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.545 0.070 174.615 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.865 0.070 179.935 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.185 0.070 185.255 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.505 0.070 190.575 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.825 0.070 195.895 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.145 0.070 201.215 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.465 0.070 206.535 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.785 0.070 211.855 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.105 0.070 217.175 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.425 0.070 222.495 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.745 0.070 227.815 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.065 0.070 233.135 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.385 0.070 238.455 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.705 0.070 243.775 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.025 0.070 249.095 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.345 0.070 254.415 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.665 0.070 259.735 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.985 0.070 265.055 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.305 0.070 270.375 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.625 0.070 275.695 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.945 0.070 281.015 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.265 0.070 286.335 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.585 0.070 291.655 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.905 0.070 296.975 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.225 0.070 302.295 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.545 0.070 307.615 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.865 0.070 312.935 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.185 0.070 318.255 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.505 0.070 323.575 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.825 0.070 328.895 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.145 0.070 334.215 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.085 0.070 337.155 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.405 0.070 342.475 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.725 0.070 347.795 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.045 0.070 353.115 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.365 0.070 358.435 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.685 0.070 363.755 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.005 0.070 369.075 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.325 0.070 374.395 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.645 0.070 379.715 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.965 0.070 385.035 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.285 0.070 390.355 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.605 0.070 395.675 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 400.925 0.070 400.995 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 406.245 0.070 406.315 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.565 0.070 411.635 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.885 0.070 416.955 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 422.205 0.070 422.275 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 427.525 0.070 427.595 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 432.845 0.070 432.915 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 438.165 0.070 438.235 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.485 0.070 443.555 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 448.805 0.070 448.875 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 454.125 0.070 454.195 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 459.445 0.070 459.515 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 464.765 0.070 464.835 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 470.085 0.070 470.155 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.405 0.070 475.475 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 480.725 0.070 480.795 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 486.045 0.070 486.115 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 491.365 0.070 491.435 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 496.685 0.070 496.755 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 502.005 0.070 502.075 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.945 0.070 505.015 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.265 0.070 510.335 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.585 0.070 515.655 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.905 0.070 520.975 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.225 0.070 526.295 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.545 0.070 531.615 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.865 0.070 536.935 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.185 0.070 542.255 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.505 0.070 547.575 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.825 0.070 552.895 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.145 0.070 558.215 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.465 0.070 563.535 ;
    END
  END addr_in[11]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.785 0.070 568.855 ;
    END
  END addr_in[12]
  PIN addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.105 0.070 574.175 ;
    END
  END addr_in[13]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.045 0.070 577.115 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.365 0.070 582.435 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.685 0.070 587.755 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 614.600 ;
      RECT 3.500 1.400 3.780 614.600 ;
      RECT 5.740 1.400 6.020 614.600 ;
      RECT 7.980 1.400 8.260 614.600 ;
      RECT 10.220 1.400 10.500 614.600 ;
      RECT 12.460 1.400 12.740 614.600 ;
      RECT 14.700 1.400 14.980 614.600 ;
      RECT 16.940 1.400 17.220 614.600 ;
      RECT 19.180 1.400 19.460 614.600 ;
      RECT 21.420 1.400 21.700 614.600 ;
      RECT 23.660 1.400 23.940 614.600 ;
      RECT 25.900 1.400 26.180 614.600 ;
      RECT 28.140 1.400 28.420 614.600 ;
      RECT 30.380 1.400 30.660 614.600 ;
      RECT 32.620 1.400 32.900 614.600 ;
      RECT 34.860 1.400 35.140 614.600 ;
      RECT 37.100 1.400 37.380 614.600 ;
      RECT 39.340 1.400 39.620 614.600 ;
      RECT 41.580 1.400 41.860 614.600 ;
      RECT 43.820 1.400 44.100 614.600 ;
      RECT 46.060 1.400 46.340 614.600 ;
      RECT 48.300 1.400 48.580 614.600 ;
      RECT 50.540 1.400 50.820 614.600 ;
      RECT 52.780 1.400 53.060 614.600 ;
      RECT 55.020 1.400 55.300 614.600 ;
      RECT 57.260 1.400 57.540 614.600 ;
      RECT 59.500 1.400 59.780 614.600 ;
      RECT 61.740 1.400 62.020 614.600 ;
      RECT 63.980 1.400 64.260 614.600 ;
      RECT 66.220 1.400 66.500 614.600 ;
      RECT 68.460 1.400 68.740 614.600 ;
      RECT 70.700 1.400 70.980 614.600 ;
      RECT 72.940 1.400 73.220 614.600 ;
      RECT 75.180 1.400 75.460 614.600 ;
      RECT 77.420 1.400 77.700 614.600 ;
      RECT 79.660 1.400 79.940 614.600 ;
      RECT 81.900 1.400 82.180 614.600 ;
      RECT 84.140 1.400 84.420 614.600 ;
      RECT 86.380 1.400 86.660 614.600 ;
      RECT 88.620 1.400 88.900 614.600 ;
      RECT 90.860 1.400 91.140 614.600 ;
      RECT 93.100 1.400 93.380 614.600 ;
      RECT 95.340 1.400 95.620 614.600 ;
      RECT 97.580 1.400 97.860 614.600 ;
      RECT 99.820 1.400 100.100 614.600 ;
      RECT 102.060 1.400 102.340 614.600 ;
      RECT 104.300 1.400 104.580 614.600 ;
      RECT 106.540 1.400 106.820 614.600 ;
      RECT 108.780 1.400 109.060 614.600 ;
      RECT 111.020 1.400 111.300 614.600 ;
      RECT 113.260 1.400 113.540 614.600 ;
      RECT 115.500 1.400 115.780 614.600 ;
      RECT 117.740 1.400 118.020 614.600 ;
      RECT 119.980 1.400 120.260 614.600 ;
      RECT 122.220 1.400 122.500 614.600 ;
      RECT 124.460 1.400 124.740 614.600 ;
      RECT 126.700 1.400 126.980 614.600 ;
      RECT 128.940 1.400 129.220 614.600 ;
      RECT 131.180 1.400 131.460 614.600 ;
      RECT 133.420 1.400 133.700 614.600 ;
      RECT 135.660 1.400 135.940 614.600 ;
      RECT 137.900 1.400 138.180 614.600 ;
      RECT 140.140 1.400 140.420 614.600 ;
      RECT 142.380 1.400 142.660 614.600 ;
      RECT 144.620 1.400 144.900 614.600 ;
      RECT 146.860 1.400 147.140 614.600 ;
      RECT 149.100 1.400 149.380 614.600 ;
      RECT 151.340 1.400 151.620 614.600 ;
      RECT 153.580 1.400 153.860 614.600 ;
      RECT 155.820 1.400 156.100 614.600 ;
      RECT 158.060 1.400 158.340 614.600 ;
      RECT 160.300 1.400 160.580 614.600 ;
      RECT 162.540 1.400 162.820 614.600 ;
      RECT 164.780 1.400 165.060 614.600 ;
      RECT 167.020 1.400 167.300 614.600 ;
      RECT 169.260 1.400 169.540 614.600 ;
      RECT 171.500 1.400 171.780 614.600 ;
      RECT 173.740 1.400 174.020 614.600 ;
      RECT 175.980 1.400 176.260 614.600 ;
      RECT 178.220 1.400 178.500 614.600 ;
      RECT 180.460 1.400 180.740 614.600 ;
      RECT 182.700 1.400 182.980 614.600 ;
      RECT 184.940 1.400 185.220 614.600 ;
      RECT 187.180 1.400 187.460 614.600 ;
      RECT 189.420 1.400 189.700 614.600 ;
      RECT 191.660 1.400 191.940 614.600 ;
      RECT 193.900 1.400 194.180 614.600 ;
      RECT 196.140 1.400 196.420 614.600 ;
      RECT 198.380 1.400 198.660 614.600 ;
      RECT 200.620 1.400 200.900 614.600 ;
      RECT 202.860 1.400 203.140 614.600 ;
      RECT 205.100 1.400 205.380 614.600 ;
      RECT 207.340 1.400 207.620 614.600 ;
      RECT 209.580 1.400 209.860 614.600 ;
      RECT 211.820 1.400 212.100 614.600 ;
      RECT 214.060 1.400 214.340 614.600 ;
      RECT 216.300 1.400 216.580 614.600 ;
      RECT 218.540 1.400 218.820 614.600 ;
      RECT 220.780 1.400 221.060 614.600 ;
      RECT 223.020 1.400 223.300 614.600 ;
      RECT 225.260 1.400 225.540 614.600 ;
      RECT 227.500 1.400 227.780 614.600 ;
      RECT 229.740 1.400 230.020 614.600 ;
      RECT 231.980 1.400 232.260 614.600 ;
      RECT 234.220 1.400 234.500 614.600 ;
      RECT 236.460 1.400 236.740 614.600 ;
      RECT 238.700 1.400 238.980 614.600 ;
      RECT 240.940 1.400 241.220 614.600 ;
      RECT 243.180 1.400 243.460 614.600 ;
      RECT 245.420 1.400 245.700 614.600 ;
      RECT 247.660 1.400 247.940 614.600 ;
      RECT 249.900 1.400 250.180 614.600 ;
      RECT 252.140 1.400 252.420 614.600 ;
      RECT 254.380 1.400 254.660 614.600 ;
      RECT 256.620 1.400 256.900 614.600 ;
      RECT 258.860 1.400 259.140 614.600 ;
      RECT 261.100 1.400 261.380 614.600 ;
      RECT 263.340 1.400 263.620 614.600 ;
      RECT 265.580 1.400 265.860 614.600 ;
      RECT 267.820 1.400 268.100 614.600 ;
      RECT 270.060 1.400 270.340 614.600 ;
      RECT 272.300 1.400 272.580 614.600 ;
      RECT 274.540 1.400 274.820 614.600 ;
      RECT 276.780 1.400 277.060 614.600 ;
      RECT 279.020 1.400 279.300 614.600 ;
      RECT 281.260 1.400 281.540 614.600 ;
      RECT 283.500 1.400 283.780 614.600 ;
      RECT 285.740 1.400 286.020 614.600 ;
      RECT 287.980 1.400 288.260 614.600 ;
      RECT 290.220 1.400 290.500 614.600 ;
      RECT 292.460 1.400 292.740 614.600 ;
      RECT 294.700 1.400 294.980 614.600 ;
      RECT 296.940 1.400 297.220 614.600 ;
      RECT 299.180 1.400 299.460 614.600 ;
      RECT 301.420 1.400 301.700 614.600 ;
      RECT 303.660 1.400 303.940 614.600 ;
      RECT 305.900 1.400 306.180 614.600 ;
      RECT 308.140 1.400 308.420 614.600 ;
      RECT 310.380 1.400 310.660 614.600 ;
      RECT 312.620 1.400 312.900 614.600 ;
      RECT 314.860 1.400 315.140 614.600 ;
      RECT 317.100 1.400 317.380 614.600 ;
      RECT 319.340 1.400 319.620 614.600 ;
      RECT 321.580 1.400 321.860 614.600 ;
      RECT 323.820 1.400 324.100 614.600 ;
      RECT 326.060 1.400 326.340 614.600 ;
      RECT 328.300 1.400 328.580 614.600 ;
      RECT 330.540 1.400 330.820 614.600 ;
      RECT 332.780 1.400 333.060 614.600 ;
      RECT 335.020 1.400 335.300 614.600 ;
      RECT 337.260 1.400 337.540 614.600 ;
      RECT 339.500 1.400 339.780 614.600 ;
      RECT 341.740 1.400 342.020 614.600 ;
      RECT 343.980 1.400 344.260 614.600 ;
      RECT 346.220 1.400 346.500 614.600 ;
      RECT 348.460 1.400 348.740 614.600 ;
      RECT 350.700 1.400 350.980 614.600 ;
      RECT 352.940 1.400 353.220 614.600 ;
      RECT 355.180 1.400 355.460 614.600 ;
      RECT 357.420 1.400 357.700 614.600 ;
      RECT 359.660 1.400 359.940 614.600 ;
      RECT 361.900 1.400 362.180 614.600 ;
      RECT 364.140 1.400 364.420 614.600 ;
      RECT 366.380 1.400 366.660 614.600 ;
      RECT 368.620 1.400 368.900 614.600 ;
      RECT 370.860 1.400 371.140 614.600 ;
      RECT 373.100 1.400 373.380 614.600 ;
      RECT 375.340 1.400 375.620 614.600 ;
      RECT 377.580 1.400 377.860 614.600 ;
      RECT 379.820 1.400 380.100 614.600 ;
      RECT 382.060 1.400 382.340 614.600 ;
      RECT 384.300 1.400 384.580 614.600 ;
      RECT 386.540 1.400 386.820 614.600 ;
      RECT 388.780 1.400 389.060 614.600 ;
      RECT 391.020 1.400 391.300 614.600 ;
      RECT 393.260 1.400 393.540 614.600 ;
      RECT 395.500 1.400 395.780 614.600 ;
      RECT 397.740 1.400 398.020 614.600 ;
      RECT 399.980 1.400 400.260 614.600 ;
      RECT 402.220 1.400 402.500 614.600 ;
      RECT 404.460 1.400 404.740 614.600 ;
      RECT 406.700 1.400 406.980 614.600 ;
      RECT 408.940 1.400 409.220 614.600 ;
      RECT 411.180 1.400 411.460 614.600 ;
      RECT 413.420 1.400 413.700 614.600 ;
      RECT 415.660 1.400 415.940 614.600 ;
      RECT 417.900 1.400 418.180 614.600 ;
      RECT 420.140 1.400 420.420 614.600 ;
      RECT 422.380 1.400 422.660 614.600 ;
      RECT 424.620 1.400 424.900 614.600 ;
      RECT 426.860 1.400 427.140 614.600 ;
      RECT 429.100 1.400 429.380 614.600 ;
      RECT 431.340 1.400 431.620 614.600 ;
      RECT 433.580 1.400 433.860 614.600 ;
      RECT 435.820 1.400 436.100 614.600 ;
      RECT 438.060 1.400 438.340 614.600 ;
      RECT 440.300 1.400 440.580 614.600 ;
      RECT 442.540 1.400 442.820 614.600 ;
      RECT 444.780 1.400 445.060 614.600 ;
      RECT 447.020 1.400 447.300 614.600 ;
      RECT 449.260 1.400 449.540 614.600 ;
      RECT 451.500 1.400 451.780 614.600 ;
      RECT 453.740 1.400 454.020 614.600 ;
      RECT 455.980 1.400 456.260 614.600 ;
      RECT 458.220 1.400 458.500 614.600 ;
      RECT 460.460 1.400 460.740 614.600 ;
      RECT 462.700 1.400 462.980 614.600 ;
      RECT 464.940 1.400 465.220 614.600 ;
      RECT 467.180 1.400 467.460 614.600 ;
      RECT 469.420 1.400 469.700 614.600 ;
      RECT 471.660 1.400 471.940 614.600 ;
      RECT 473.900 1.400 474.180 614.600 ;
      RECT 476.140 1.400 476.420 614.600 ;
      RECT 478.380 1.400 478.660 614.600 ;
      RECT 480.620 1.400 480.900 614.600 ;
      RECT 482.860 1.400 483.140 614.600 ;
      RECT 485.100 1.400 485.380 614.600 ;
      RECT 487.340 1.400 487.620 614.600 ;
      RECT 489.580 1.400 489.860 614.600 ;
      RECT 491.820 1.400 492.100 614.600 ;
      RECT 494.060 1.400 494.340 614.600 ;
      RECT 496.300 1.400 496.580 614.600 ;
      RECT 498.540 1.400 498.820 614.600 ;
      RECT 500.780 1.400 501.060 614.600 ;
      RECT 503.020 1.400 503.300 614.600 ;
      RECT 505.260 1.400 505.540 614.600 ;
      RECT 507.500 1.400 507.780 614.600 ;
      RECT 509.740 1.400 510.020 614.600 ;
      RECT 511.980 1.400 512.260 614.600 ;
      RECT 514.220 1.400 514.500 614.600 ;
      RECT 516.460 1.400 516.740 614.600 ;
      RECT 518.700 1.400 518.980 614.600 ;
      RECT 520.940 1.400 521.220 614.600 ;
      RECT 523.180 1.400 523.460 614.600 ;
      RECT 525.420 1.400 525.700 614.600 ;
      RECT 527.660 1.400 527.940 614.600 ;
      RECT 529.900 1.400 530.180 614.600 ;
      RECT 532.140 1.400 532.420 614.600 ;
      RECT 534.380 1.400 534.660 614.600 ;
      RECT 536.620 1.400 536.900 614.600 ;
      RECT 538.860 1.400 539.140 614.600 ;
      RECT 541.100 1.400 541.380 614.600 ;
      RECT 543.340 1.400 543.620 614.600 ;
      RECT 545.580 1.400 545.860 614.600 ;
      RECT 547.820 1.400 548.100 614.600 ;
      RECT 550.060 1.400 550.340 614.600 ;
      RECT 552.300 1.400 552.580 614.600 ;
      RECT 554.540 1.400 554.820 614.600 ;
      RECT 556.780 1.400 557.060 614.600 ;
      RECT 559.020 1.400 559.300 614.600 ;
      RECT 561.260 1.400 561.540 614.600 ;
      RECT 563.500 1.400 563.780 614.600 ;
      RECT 565.740 1.400 566.020 614.600 ;
      RECT 567.980 1.400 568.260 614.600 ;
      RECT 570.220 1.400 570.500 614.600 ;
      RECT 572.460 1.400 572.740 614.600 ;
      RECT 574.700 1.400 574.980 614.600 ;
      RECT 576.940 1.400 577.220 614.600 ;
      RECT 579.180 1.400 579.460 614.600 ;
      RECT 581.420 1.400 581.700 614.600 ;
      RECT 583.660 1.400 583.940 614.600 ;
      RECT 585.900 1.400 586.180 614.600 ;
      RECT 588.140 1.400 588.420 614.600 ;
      RECT 590.380 1.400 590.660 614.600 ;
      RECT 592.620 1.400 592.900 614.600 ;
      RECT 594.860 1.400 595.140 614.600 ;
      RECT 597.100 1.400 597.380 614.600 ;
      RECT 599.340 1.400 599.620 614.600 ;
      RECT 601.580 1.400 601.860 614.600 ;
      RECT 603.820 1.400 604.100 614.600 ;
      RECT 606.060 1.400 606.340 614.600 ;
      RECT 608.300 1.400 608.580 614.600 ;
      RECT 610.540 1.400 610.820 614.600 ;
      RECT 612.780 1.400 613.060 614.600 ;
      RECT 615.020 1.400 615.300 614.600 ;
      RECT 617.260 1.400 617.540 614.600 ;
      RECT 619.500 1.400 619.780 614.600 ;
      RECT 621.740 1.400 622.020 614.600 ;
      RECT 623.980 1.400 624.260 614.600 ;
      RECT 626.220 1.400 626.500 614.600 ;
      RECT 628.460 1.400 628.740 614.600 ;
      RECT 630.700 1.400 630.980 614.600 ;
      RECT 632.940 1.400 633.220 614.600 ;
      RECT 635.180 1.400 635.460 614.600 ;
      RECT 637.420 1.400 637.700 614.600 ;
      RECT 639.660 1.400 639.940 614.600 ;
      RECT 641.900 1.400 642.180 614.600 ;
      RECT 644.140 1.400 644.420 614.600 ;
      RECT 646.380 1.400 646.660 614.600 ;
      RECT 648.620 1.400 648.900 614.600 ;
      RECT 650.860 1.400 651.140 614.600 ;
      RECT 653.100 1.400 653.380 614.600 ;
      RECT 655.340 1.400 655.620 614.600 ;
      RECT 657.580 1.400 657.860 614.600 ;
      RECT 659.820 1.400 660.100 614.600 ;
      RECT 662.060 1.400 662.340 614.600 ;
      RECT 664.300 1.400 664.580 614.600 ;
      RECT 666.540 1.400 666.820 614.600 ;
      RECT 668.780 1.400 669.060 614.600 ;
      RECT 671.020 1.400 671.300 614.600 ;
      RECT 673.260 1.400 673.540 614.600 ;
      RECT 675.500 1.400 675.780 614.600 ;
      RECT 677.740 1.400 678.020 614.600 ;
      RECT 679.980 1.400 680.260 614.600 ;
      RECT 682.220 1.400 682.500 614.600 ;
      RECT 684.460 1.400 684.740 614.600 ;
      RECT 686.700 1.400 686.980 614.600 ;
      RECT 688.940 1.400 689.220 614.600 ;
      RECT 691.180 1.400 691.460 614.600 ;
      RECT 693.420 1.400 693.700 614.600 ;
      RECT 695.660 1.400 695.940 614.600 ;
      RECT 697.900 1.400 698.180 614.600 ;
      RECT 700.140 1.400 700.420 614.600 ;
      RECT 702.380 1.400 702.660 614.600 ;
      RECT 704.620 1.400 704.900 614.600 ;
      RECT 706.860 1.400 707.140 614.600 ;
      RECT 709.100 1.400 709.380 614.600 ;
      RECT 711.340 1.400 711.620 614.600 ;
      RECT 713.580 1.400 713.860 614.600 ;
      RECT 715.820 1.400 716.100 614.600 ;
      RECT 718.060 1.400 718.340 614.600 ;
      RECT 720.300 1.400 720.580 614.600 ;
      RECT 722.540 1.400 722.820 614.600 ;
      RECT 724.780 1.400 725.060 614.600 ;
      RECT 727.020 1.400 727.300 614.600 ;
      RECT 729.260 1.400 729.540 614.600 ;
      RECT 731.500 1.400 731.780 614.600 ;
      RECT 733.740 1.400 734.020 614.600 ;
      RECT 735.980 1.400 736.260 614.600 ;
      RECT 738.220 1.400 738.500 614.600 ;
      RECT 740.460 1.400 740.740 614.600 ;
      RECT 742.700 1.400 742.980 614.600 ;
      RECT 744.940 1.400 745.220 614.600 ;
      RECT 747.180 1.400 747.460 614.600 ;
      RECT 749.420 1.400 749.700 614.600 ;
      RECT 751.660 1.400 751.940 614.600 ;
      RECT 753.900 1.400 754.180 614.600 ;
      RECT 756.140 1.400 756.420 614.600 ;
      RECT 758.380 1.400 758.660 614.600 ;
      RECT 760.620 1.400 760.900 614.600 ;
      RECT 762.860 1.400 763.140 614.600 ;
      RECT 765.100 1.400 765.380 614.600 ;
      RECT 767.340 1.400 767.620 614.600 ;
      RECT 769.580 1.400 769.860 614.600 ;
      RECT 771.820 1.400 772.100 614.600 ;
      RECT 774.060 1.400 774.340 614.600 ;
      RECT 776.300 1.400 776.580 614.600 ;
      RECT 778.540 1.400 778.820 614.600 ;
      RECT 780.780 1.400 781.060 614.600 ;
      RECT 783.020 1.400 783.300 614.600 ;
      RECT 785.260 1.400 785.540 614.600 ;
      RECT 787.500 1.400 787.780 614.600 ;
      RECT 789.740 1.400 790.020 614.600 ;
      RECT 791.980 1.400 792.260 614.600 ;
      RECT 794.220 1.400 794.500 614.600 ;
      RECT 796.460 1.400 796.740 614.600 ;
      RECT 798.700 1.400 798.980 614.600 ;
      RECT 800.940 1.400 801.220 614.600 ;
      RECT 803.180 1.400 803.460 614.600 ;
      RECT 805.420 1.400 805.700 614.600 ;
      RECT 807.660 1.400 807.940 614.600 ;
      RECT 809.900 1.400 810.180 614.600 ;
      RECT 812.140 1.400 812.420 614.600 ;
      RECT 814.380 1.400 814.660 614.600 ;
      RECT 816.620 1.400 816.900 614.600 ;
      RECT 818.860 1.400 819.140 614.600 ;
      RECT 821.100 1.400 821.380 614.600 ;
      RECT 823.340 1.400 823.620 614.600 ;
      RECT 825.580 1.400 825.860 614.600 ;
      RECT 827.820 1.400 828.100 614.600 ;
      RECT 830.060 1.400 830.340 614.600 ;
      RECT 832.300 1.400 832.580 614.600 ;
      RECT 834.540 1.400 834.820 614.600 ;
      RECT 836.780 1.400 837.060 614.600 ;
      RECT 839.020 1.400 839.300 614.600 ;
      RECT 841.260 1.400 841.540 614.600 ;
      RECT 843.500 1.400 843.780 614.600 ;
      RECT 845.740 1.400 846.020 614.600 ;
      RECT 847.980 1.400 848.260 614.600 ;
      RECT 850.220 1.400 850.500 614.600 ;
      RECT 852.460 1.400 852.740 614.600 ;
      RECT 854.700 1.400 854.980 614.600 ;
      RECT 856.940 1.400 857.220 614.600 ;
      RECT 859.180 1.400 859.460 614.600 ;
      RECT 861.420 1.400 861.700 614.600 ;
      RECT 863.660 1.400 863.940 614.600 ;
      RECT 865.900 1.400 866.180 614.600 ;
      RECT 868.140 1.400 868.420 614.600 ;
      RECT 870.380 1.400 870.660 614.600 ;
      RECT 872.620 1.400 872.900 614.600 ;
      RECT 874.860 1.400 875.140 614.600 ;
      RECT 877.100 1.400 877.380 614.600 ;
      RECT 879.340 1.400 879.620 614.600 ;
      RECT 881.580 1.400 881.860 614.600 ;
      RECT 883.820 1.400 884.100 614.600 ;
      RECT 886.060 1.400 886.340 614.600 ;
      RECT 888.300 1.400 888.580 614.600 ;
      RECT 890.540 1.400 890.820 614.600 ;
      RECT 892.780 1.400 893.060 614.600 ;
      RECT 895.020 1.400 895.300 614.600 ;
      RECT 897.260 1.400 897.540 614.600 ;
      RECT 899.500 1.400 899.780 614.600 ;
      RECT 901.740 1.400 902.020 614.600 ;
      RECT 903.980 1.400 904.260 614.600 ;
      RECT 906.220 1.400 906.500 614.600 ;
      RECT 908.460 1.400 908.740 614.600 ;
      RECT 910.700 1.400 910.980 614.600 ;
      RECT 912.940 1.400 913.220 614.600 ;
      RECT 915.180 1.400 915.460 614.600 ;
      RECT 917.420 1.400 917.700 614.600 ;
      RECT 919.660 1.400 919.940 614.600 ;
      RECT 921.900 1.400 922.180 614.600 ;
      RECT 924.140 1.400 924.420 614.600 ;
      RECT 926.380 1.400 926.660 614.600 ;
      RECT 928.620 1.400 928.900 614.600 ;
      RECT 930.860 1.400 931.140 614.600 ;
      RECT 933.100 1.400 933.380 614.600 ;
      RECT 935.340 1.400 935.620 614.600 ;
      RECT 937.580 1.400 937.860 614.600 ;
      RECT 939.820 1.400 940.100 614.600 ;
      RECT 942.060 1.400 942.340 614.600 ;
      RECT 944.300 1.400 944.580 614.600 ;
      RECT 946.540 1.400 946.820 614.600 ;
      RECT 948.780 1.400 949.060 614.600 ;
      RECT 951.020 1.400 951.300 614.600 ;
      RECT 953.260 1.400 953.540 614.600 ;
      RECT 955.500 1.400 955.780 614.600 ;
      RECT 957.740 1.400 958.020 614.600 ;
      RECT 959.980 1.400 960.260 614.600 ;
      RECT 962.220 1.400 962.500 614.600 ;
      RECT 964.460 1.400 964.740 614.600 ;
      RECT 966.700 1.400 966.980 614.600 ;
      RECT 968.940 1.400 969.220 614.600 ;
      RECT 971.180 1.400 971.460 614.600 ;
      RECT 973.420 1.400 973.700 614.600 ;
      RECT 975.660 1.400 975.940 614.600 ;
      RECT 977.900 1.400 978.180 614.600 ;
      RECT 980.140 1.400 980.420 614.600 ;
      RECT 982.380 1.400 982.660 614.600 ;
      RECT 984.620 1.400 984.900 614.600 ;
      RECT 986.860 1.400 987.140 614.600 ;
      RECT 989.100 1.400 989.380 614.600 ;
      RECT 991.340 1.400 991.620 614.600 ;
      RECT 993.580 1.400 993.860 614.600 ;
      RECT 995.820 1.400 996.100 614.600 ;
      RECT 998.060 1.400 998.340 614.600 ;
      RECT 1000.300 1.400 1000.580 614.600 ;
      RECT 1002.540 1.400 1002.820 614.600 ;
      RECT 1004.780 1.400 1005.060 614.600 ;
      RECT 1007.020 1.400 1007.300 614.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 614.600 ;
      RECT 4.620 1.400 4.900 614.600 ;
      RECT 6.860 1.400 7.140 614.600 ;
      RECT 9.100 1.400 9.380 614.600 ;
      RECT 11.340 1.400 11.620 614.600 ;
      RECT 13.580 1.400 13.860 614.600 ;
      RECT 15.820 1.400 16.100 614.600 ;
      RECT 18.060 1.400 18.340 614.600 ;
      RECT 20.300 1.400 20.580 614.600 ;
      RECT 22.540 1.400 22.820 614.600 ;
      RECT 24.780 1.400 25.060 614.600 ;
      RECT 27.020 1.400 27.300 614.600 ;
      RECT 29.260 1.400 29.540 614.600 ;
      RECT 31.500 1.400 31.780 614.600 ;
      RECT 33.740 1.400 34.020 614.600 ;
      RECT 35.980 1.400 36.260 614.600 ;
      RECT 38.220 1.400 38.500 614.600 ;
      RECT 40.460 1.400 40.740 614.600 ;
      RECT 42.700 1.400 42.980 614.600 ;
      RECT 44.940 1.400 45.220 614.600 ;
      RECT 47.180 1.400 47.460 614.600 ;
      RECT 49.420 1.400 49.700 614.600 ;
      RECT 51.660 1.400 51.940 614.600 ;
      RECT 53.900 1.400 54.180 614.600 ;
      RECT 56.140 1.400 56.420 614.600 ;
      RECT 58.380 1.400 58.660 614.600 ;
      RECT 60.620 1.400 60.900 614.600 ;
      RECT 62.860 1.400 63.140 614.600 ;
      RECT 65.100 1.400 65.380 614.600 ;
      RECT 67.340 1.400 67.620 614.600 ;
      RECT 69.580 1.400 69.860 614.600 ;
      RECT 71.820 1.400 72.100 614.600 ;
      RECT 74.060 1.400 74.340 614.600 ;
      RECT 76.300 1.400 76.580 614.600 ;
      RECT 78.540 1.400 78.820 614.600 ;
      RECT 80.780 1.400 81.060 614.600 ;
      RECT 83.020 1.400 83.300 614.600 ;
      RECT 85.260 1.400 85.540 614.600 ;
      RECT 87.500 1.400 87.780 614.600 ;
      RECT 89.740 1.400 90.020 614.600 ;
      RECT 91.980 1.400 92.260 614.600 ;
      RECT 94.220 1.400 94.500 614.600 ;
      RECT 96.460 1.400 96.740 614.600 ;
      RECT 98.700 1.400 98.980 614.600 ;
      RECT 100.940 1.400 101.220 614.600 ;
      RECT 103.180 1.400 103.460 614.600 ;
      RECT 105.420 1.400 105.700 614.600 ;
      RECT 107.660 1.400 107.940 614.600 ;
      RECT 109.900 1.400 110.180 614.600 ;
      RECT 112.140 1.400 112.420 614.600 ;
      RECT 114.380 1.400 114.660 614.600 ;
      RECT 116.620 1.400 116.900 614.600 ;
      RECT 118.860 1.400 119.140 614.600 ;
      RECT 121.100 1.400 121.380 614.600 ;
      RECT 123.340 1.400 123.620 614.600 ;
      RECT 125.580 1.400 125.860 614.600 ;
      RECT 127.820 1.400 128.100 614.600 ;
      RECT 130.060 1.400 130.340 614.600 ;
      RECT 132.300 1.400 132.580 614.600 ;
      RECT 134.540 1.400 134.820 614.600 ;
      RECT 136.780 1.400 137.060 614.600 ;
      RECT 139.020 1.400 139.300 614.600 ;
      RECT 141.260 1.400 141.540 614.600 ;
      RECT 143.500 1.400 143.780 614.600 ;
      RECT 145.740 1.400 146.020 614.600 ;
      RECT 147.980 1.400 148.260 614.600 ;
      RECT 150.220 1.400 150.500 614.600 ;
      RECT 152.460 1.400 152.740 614.600 ;
      RECT 154.700 1.400 154.980 614.600 ;
      RECT 156.940 1.400 157.220 614.600 ;
      RECT 159.180 1.400 159.460 614.600 ;
      RECT 161.420 1.400 161.700 614.600 ;
      RECT 163.660 1.400 163.940 614.600 ;
      RECT 165.900 1.400 166.180 614.600 ;
      RECT 168.140 1.400 168.420 614.600 ;
      RECT 170.380 1.400 170.660 614.600 ;
      RECT 172.620 1.400 172.900 614.600 ;
      RECT 174.860 1.400 175.140 614.600 ;
      RECT 177.100 1.400 177.380 614.600 ;
      RECT 179.340 1.400 179.620 614.600 ;
      RECT 181.580 1.400 181.860 614.600 ;
      RECT 183.820 1.400 184.100 614.600 ;
      RECT 186.060 1.400 186.340 614.600 ;
      RECT 188.300 1.400 188.580 614.600 ;
      RECT 190.540 1.400 190.820 614.600 ;
      RECT 192.780 1.400 193.060 614.600 ;
      RECT 195.020 1.400 195.300 614.600 ;
      RECT 197.260 1.400 197.540 614.600 ;
      RECT 199.500 1.400 199.780 614.600 ;
      RECT 201.740 1.400 202.020 614.600 ;
      RECT 203.980 1.400 204.260 614.600 ;
      RECT 206.220 1.400 206.500 614.600 ;
      RECT 208.460 1.400 208.740 614.600 ;
      RECT 210.700 1.400 210.980 614.600 ;
      RECT 212.940 1.400 213.220 614.600 ;
      RECT 215.180 1.400 215.460 614.600 ;
      RECT 217.420 1.400 217.700 614.600 ;
      RECT 219.660 1.400 219.940 614.600 ;
      RECT 221.900 1.400 222.180 614.600 ;
      RECT 224.140 1.400 224.420 614.600 ;
      RECT 226.380 1.400 226.660 614.600 ;
      RECT 228.620 1.400 228.900 614.600 ;
      RECT 230.860 1.400 231.140 614.600 ;
      RECT 233.100 1.400 233.380 614.600 ;
      RECT 235.340 1.400 235.620 614.600 ;
      RECT 237.580 1.400 237.860 614.600 ;
      RECT 239.820 1.400 240.100 614.600 ;
      RECT 242.060 1.400 242.340 614.600 ;
      RECT 244.300 1.400 244.580 614.600 ;
      RECT 246.540 1.400 246.820 614.600 ;
      RECT 248.780 1.400 249.060 614.600 ;
      RECT 251.020 1.400 251.300 614.600 ;
      RECT 253.260 1.400 253.540 614.600 ;
      RECT 255.500 1.400 255.780 614.600 ;
      RECT 257.740 1.400 258.020 614.600 ;
      RECT 259.980 1.400 260.260 614.600 ;
      RECT 262.220 1.400 262.500 614.600 ;
      RECT 264.460 1.400 264.740 614.600 ;
      RECT 266.700 1.400 266.980 614.600 ;
      RECT 268.940 1.400 269.220 614.600 ;
      RECT 271.180 1.400 271.460 614.600 ;
      RECT 273.420 1.400 273.700 614.600 ;
      RECT 275.660 1.400 275.940 614.600 ;
      RECT 277.900 1.400 278.180 614.600 ;
      RECT 280.140 1.400 280.420 614.600 ;
      RECT 282.380 1.400 282.660 614.600 ;
      RECT 284.620 1.400 284.900 614.600 ;
      RECT 286.860 1.400 287.140 614.600 ;
      RECT 289.100 1.400 289.380 614.600 ;
      RECT 291.340 1.400 291.620 614.600 ;
      RECT 293.580 1.400 293.860 614.600 ;
      RECT 295.820 1.400 296.100 614.600 ;
      RECT 298.060 1.400 298.340 614.600 ;
      RECT 300.300 1.400 300.580 614.600 ;
      RECT 302.540 1.400 302.820 614.600 ;
      RECT 304.780 1.400 305.060 614.600 ;
      RECT 307.020 1.400 307.300 614.600 ;
      RECT 309.260 1.400 309.540 614.600 ;
      RECT 311.500 1.400 311.780 614.600 ;
      RECT 313.740 1.400 314.020 614.600 ;
      RECT 315.980 1.400 316.260 614.600 ;
      RECT 318.220 1.400 318.500 614.600 ;
      RECT 320.460 1.400 320.740 614.600 ;
      RECT 322.700 1.400 322.980 614.600 ;
      RECT 324.940 1.400 325.220 614.600 ;
      RECT 327.180 1.400 327.460 614.600 ;
      RECT 329.420 1.400 329.700 614.600 ;
      RECT 331.660 1.400 331.940 614.600 ;
      RECT 333.900 1.400 334.180 614.600 ;
      RECT 336.140 1.400 336.420 614.600 ;
      RECT 338.380 1.400 338.660 614.600 ;
      RECT 340.620 1.400 340.900 614.600 ;
      RECT 342.860 1.400 343.140 614.600 ;
      RECT 345.100 1.400 345.380 614.600 ;
      RECT 347.340 1.400 347.620 614.600 ;
      RECT 349.580 1.400 349.860 614.600 ;
      RECT 351.820 1.400 352.100 614.600 ;
      RECT 354.060 1.400 354.340 614.600 ;
      RECT 356.300 1.400 356.580 614.600 ;
      RECT 358.540 1.400 358.820 614.600 ;
      RECT 360.780 1.400 361.060 614.600 ;
      RECT 363.020 1.400 363.300 614.600 ;
      RECT 365.260 1.400 365.540 614.600 ;
      RECT 367.500 1.400 367.780 614.600 ;
      RECT 369.740 1.400 370.020 614.600 ;
      RECT 371.980 1.400 372.260 614.600 ;
      RECT 374.220 1.400 374.500 614.600 ;
      RECT 376.460 1.400 376.740 614.600 ;
      RECT 378.700 1.400 378.980 614.600 ;
      RECT 380.940 1.400 381.220 614.600 ;
      RECT 383.180 1.400 383.460 614.600 ;
      RECT 385.420 1.400 385.700 614.600 ;
      RECT 387.660 1.400 387.940 614.600 ;
      RECT 389.900 1.400 390.180 614.600 ;
      RECT 392.140 1.400 392.420 614.600 ;
      RECT 394.380 1.400 394.660 614.600 ;
      RECT 396.620 1.400 396.900 614.600 ;
      RECT 398.860 1.400 399.140 614.600 ;
      RECT 401.100 1.400 401.380 614.600 ;
      RECT 403.340 1.400 403.620 614.600 ;
      RECT 405.580 1.400 405.860 614.600 ;
      RECT 407.820 1.400 408.100 614.600 ;
      RECT 410.060 1.400 410.340 614.600 ;
      RECT 412.300 1.400 412.580 614.600 ;
      RECT 414.540 1.400 414.820 614.600 ;
      RECT 416.780 1.400 417.060 614.600 ;
      RECT 419.020 1.400 419.300 614.600 ;
      RECT 421.260 1.400 421.540 614.600 ;
      RECT 423.500 1.400 423.780 614.600 ;
      RECT 425.740 1.400 426.020 614.600 ;
      RECT 427.980 1.400 428.260 614.600 ;
      RECT 430.220 1.400 430.500 614.600 ;
      RECT 432.460 1.400 432.740 614.600 ;
      RECT 434.700 1.400 434.980 614.600 ;
      RECT 436.940 1.400 437.220 614.600 ;
      RECT 439.180 1.400 439.460 614.600 ;
      RECT 441.420 1.400 441.700 614.600 ;
      RECT 443.660 1.400 443.940 614.600 ;
      RECT 445.900 1.400 446.180 614.600 ;
      RECT 448.140 1.400 448.420 614.600 ;
      RECT 450.380 1.400 450.660 614.600 ;
      RECT 452.620 1.400 452.900 614.600 ;
      RECT 454.860 1.400 455.140 614.600 ;
      RECT 457.100 1.400 457.380 614.600 ;
      RECT 459.340 1.400 459.620 614.600 ;
      RECT 461.580 1.400 461.860 614.600 ;
      RECT 463.820 1.400 464.100 614.600 ;
      RECT 466.060 1.400 466.340 614.600 ;
      RECT 468.300 1.400 468.580 614.600 ;
      RECT 470.540 1.400 470.820 614.600 ;
      RECT 472.780 1.400 473.060 614.600 ;
      RECT 475.020 1.400 475.300 614.600 ;
      RECT 477.260 1.400 477.540 614.600 ;
      RECT 479.500 1.400 479.780 614.600 ;
      RECT 481.740 1.400 482.020 614.600 ;
      RECT 483.980 1.400 484.260 614.600 ;
      RECT 486.220 1.400 486.500 614.600 ;
      RECT 488.460 1.400 488.740 614.600 ;
      RECT 490.700 1.400 490.980 614.600 ;
      RECT 492.940 1.400 493.220 614.600 ;
      RECT 495.180 1.400 495.460 614.600 ;
      RECT 497.420 1.400 497.700 614.600 ;
      RECT 499.660 1.400 499.940 614.600 ;
      RECT 501.900 1.400 502.180 614.600 ;
      RECT 504.140 1.400 504.420 614.600 ;
      RECT 506.380 1.400 506.660 614.600 ;
      RECT 508.620 1.400 508.900 614.600 ;
      RECT 510.860 1.400 511.140 614.600 ;
      RECT 513.100 1.400 513.380 614.600 ;
      RECT 515.340 1.400 515.620 614.600 ;
      RECT 517.580 1.400 517.860 614.600 ;
      RECT 519.820 1.400 520.100 614.600 ;
      RECT 522.060 1.400 522.340 614.600 ;
      RECT 524.300 1.400 524.580 614.600 ;
      RECT 526.540 1.400 526.820 614.600 ;
      RECT 528.780 1.400 529.060 614.600 ;
      RECT 531.020 1.400 531.300 614.600 ;
      RECT 533.260 1.400 533.540 614.600 ;
      RECT 535.500 1.400 535.780 614.600 ;
      RECT 537.740 1.400 538.020 614.600 ;
      RECT 539.980 1.400 540.260 614.600 ;
      RECT 542.220 1.400 542.500 614.600 ;
      RECT 544.460 1.400 544.740 614.600 ;
      RECT 546.700 1.400 546.980 614.600 ;
      RECT 548.940 1.400 549.220 614.600 ;
      RECT 551.180 1.400 551.460 614.600 ;
      RECT 553.420 1.400 553.700 614.600 ;
      RECT 555.660 1.400 555.940 614.600 ;
      RECT 557.900 1.400 558.180 614.600 ;
      RECT 560.140 1.400 560.420 614.600 ;
      RECT 562.380 1.400 562.660 614.600 ;
      RECT 564.620 1.400 564.900 614.600 ;
      RECT 566.860 1.400 567.140 614.600 ;
      RECT 569.100 1.400 569.380 614.600 ;
      RECT 571.340 1.400 571.620 614.600 ;
      RECT 573.580 1.400 573.860 614.600 ;
      RECT 575.820 1.400 576.100 614.600 ;
      RECT 578.060 1.400 578.340 614.600 ;
      RECT 580.300 1.400 580.580 614.600 ;
      RECT 582.540 1.400 582.820 614.600 ;
      RECT 584.780 1.400 585.060 614.600 ;
      RECT 587.020 1.400 587.300 614.600 ;
      RECT 589.260 1.400 589.540 614.600 ;
      RECT 591.500 1.400 591.780 614.600 ;
      RECT 593.740 1.400 594.020 614.600 ;
      RECT 595.980 1.400 596.260 614.600 ;
      RECT 598.220 1.400 598.500 614.600 ;
      RECT 600.460 1.400 600.740 614.600 ;
      RECT 602.700 1.400 602.980 614.600 ;
      RECT 604.940 1.400 605.220 614.600 ;
      RECT 607.180 1.400 607.460 614.600 ;
      RECT 609.420 1.400 609.700 614.600 ;
      RECT 611.660 1.400 611.940 614.600 ;
      RECT 613.900 1.400 614.180 614.600 ;
      RECT 616.140 1.400 616.420 614.600 ;
      RECT 618.380 1.400 618.660 614.600 ;
      RECT 620.620 1.400 620.900 614.600 ;
      RECT 622.860 1.400 623.140 614.600 ;
      RECT 625.100 1.400 625.380 614.600 ;
      RECT 627.340 1.400 627.620 614.600 ;
      RECT 629.580 1.400 629.860 614.600 ;
      RECT 631.820 1.400 632.100 614.600 ;
      RECT 634.060 1.400 634.340 614.600 ;
      RECT 636.300 1.400 636.580 614.600 ;
      RECT 638.540 1.400 638.820 614.600 ;
      RECT 640.780 1.400 641.060 614.600 ;
      RECT 643.020 1.400 643.300 614.600 ;
      RECT 645.260 1.400 645.540 614.600 ;
      RECT 647.500 1.400 647.780 614.600 ;
      RECT 649.740 1.400 650.020 614.600 ;
      RECT 651.980 1.400 652.260 614.600 ;
      RECT 654.220 1.400 654.500 614.600 ;
      RECT 656.460 1.400 656.740 614.600 ;
      RECT 658.700 1.400 658.980 614.600 ;
      RECT 660.940 1.400 661.220 614.600 ;
      RECT 663.180 1.400 663.460 614.600 ;
      RECT 665.420 1.400 665.700 614.600 ;
      RECT 667.660 1.400 667.940 614.600 ;
      RECT 669.900 1.400 670.180 614.600 ;
      RECT 672.140 1.400 672.420 614.600 ;
      RECT 674.380 1.400 674.660 614.600 ;
      RECT 676.620 1.400 676.900 614.600 ;
      RECT 678.860 1.400 679.140 614.600 ;
      RECT 681.100 1.400 681.380 614.600 ;
      RECT 683.340 1.400 683.620 614.600 ;
      RECT 685.580 1.400 685.860 614.600 ;
      RECT 687.820 1.400 688.100 614.600 ;
      RECT 690.060 1.400 690.340 614.600 ;
      RECT 692.300 1.400 692.580 614.600 ;
      RECT 694.540 1.400 694.820 614.600 ;
      RECT 696.780 1.400 697.060 614.600 ;
      RECT 699.020 1.400 699.300 614.600 ;
      RECT 701.260 1.400 701.540 614.600 ;
      RECT 703.500 1.400 703.780 614.600 ;
      RECT 705.740 1.400 706.020 614.600 ;
      RECT 707.980 1.400 708.260 614.600 ;
      RECT 710.220 1.400 710.500 614.600 ;
      RECT 712.460 1.400 712.740 614.600 ;
      RECT 714.700 1.400 714.980 614.600 ;
      RECT 716.940 1.400 717.220 614.600 ;
      RECT 719.180 1.400 719.460 614.600 ;
      RECT 721.420 1.400 721.700 614.600 ;
      RECT 723.660 1.400 723.940 614.600 ;
      RECT 725.900 1.400 726.180 614.600 ;
      RECT 728.140 1.400 728.420 614.600 ;
      RECT 730.380 1.400 730.660 614.600 ;
      RECT 732.620 1.400 732.900 614.600 ;
      RECT 734.860 1.400 735.140 614.600 ;
      RECT 737.100 1.400 737.380 614.600 ;
      RECT 739.340 1.400 739.620 614.600 ;
      RECT 741.580 1.400 741.860 614.600 ;
      RECT 743.820 1.400 744.100 614.600 ;
      RECT 746.060 1.400 746.340 614.600 ;
      RECT 748.300 1.400 748.580 614.600 ;
      RECT 750.540 1.400 750.820 614.600 ;
      RECT 752.780 1.400 753.060 614.600 ;
      RECT 755.020 1.400 755.300 614.600 ;
      RECT 757.260 1.400 757.540 614.600 ;
      RECT 759.500 1.400 759.780 614.600 ;
      RECT 761.740 1.400 762.020 614.600 ;
      RECT 763.980 1.400 764.260 614.600 ;
      RECT 766.220 1.400 766.500 614.600 ;
      RECT 768.460 1.400 768.740 614.600 ;
      RECT 770.700 1.400 770.980 614.600 ;
      RECT 772.940 1.400 773.220 614.600 ;
      RECT 775.180 1.400 775.460 614.600 ;
      RECT 777.420 1.400 777.700 614.600 ;
      RECT 779.660 1.400 779.940 614.600 ;
      RECT 781.900 1.400 782.180 614.600 ;
      RECT 784.140 1.400 784.420 614.600 ;
      RECT 786.380 1.400 786.660 614.600 ;
      RECT 788.620 1.400 788.900 614.600 ;
      RECT 790.860 1.400 791.140 614.600 ;
      RECT 793.100 1.400 793.380 614.600 ;
      RECT 795.340 1.400 795.620 614.600 ;
      RECT 797.580 1.400 797.860 614.600 ;
      RECT 799.820 1.400 800.100 614.600 ;
      RECT 802.060 1.400 802.340 614.600 ;
      RECT 804.300 1.400 804.580 614.600 ;
      RECT 806.540 1.400 806.820 614.600 ;
      RECT 808.780 1.400 809.060 614.600 ;
      RECT 811.020 1.400 811.300 614.600 ;
      RECT 813.260 1.400 813.540 614.600 ;
      RECT 815.500 1.400 815.780 614.600 ;
      RECT 817.740 1.400 818.020 614.600 ;
      RECT 819.980 1.400 820.260 614.600 ;
      RECT 822.220 1.400 822.500 614.600 ;
      RECT 824.460 1.400 824.740 614.600 ;
      RECT 826.700 1.400 826.980 614.600 ;
      RECT 828.940 1.400 829.220 614.600 ;
      RECT 831.180 1.400 831.460 614.600 ;
      RECT 833.420 1.400 833.700 614.600 ;
      RECT 835.660 1.400 835.940 614.600 ;
      RECT 837.900 1.400 838.180 614.600 ;
      RECT 840.140 1.400 840.420 614.600 ;
      RECT 842.380 1.400 842.660 614.600 ;
      RECT 844.620 1.400 844.900 614.600 ;
      RECT 846.860 1.400 847.140 614.600 ;
      RECT 849.100 1.400 849.380 614.600 ;
      RECT 851.340 1.400 851.620 614.600 ;
      RECT 853.580 1.400 853.860 614.600 ;
      RECT 855.820 1.400 856.100 614.600 ;
      RECT 858.060 1.400 858.340 614.600 ;
      RECT 860.300 1.400 860.580 614.600 ;
      RECT 862.540 1.400 862.820 614.600 ;
      RECT 864.780 1.400 865.060 614.600 ;
      RECT 867.020 1.400 867.300 614.600 ;
      RECT 869.260 1.400 869.540 614.600 ;
      RECT 871.500 1.400 871.780 614.600 ;
      RECT 873.740 1.400 874.020 614.600 ;
      RECT 875.980 1.400 876.260 614.600 ;
      RECT 878.220 1.400 878.500 614.600 ;
      RECT 880.460 1.400 880.740 614.600 ;
      RECT 882.700 1.400 882.980 614.600 ;
      RECT 884.940 1.400 885.220 614.600 ;
      RECT 887.180 1.400 887.460 614.600 ;
      RECT 889.420 1.400 889.700 614.600 ;
      RECT 891.660 1.400 891.940 614.600 ;
      RECT 893.900 1.400 894.180 614.600 ;
      RECT 896.140 1.400 896.420 614.600 ;
      RECT 898.380 1.400 898.660 614.600 ;
      RECT 900.620 1.400 900.900 614.600 ;
      RECT 902.860 1.400 903.140 614.600 ;
      RECT 905.100 1.400 905.380 614.600 ;
      RECT 907.340 1.400 907.620 614.600 ;
      RECT 909.580 1.400 909.860 614.600 ;
      RECT 911.820 1.400 912.100 614.600 ;
      RECT 914.060 1.400 914.340 614.600 ;
      RECT 916.300 1.400 916.580 614.600 ;
      RECT 918.540 1.400 918.820 614.600 ;
      RECT 920.780 1.400 921.060 614.600 ;
      RECT 923.020 1.400 923.300 614.600 ;
      RECT 925.260 1.400 925.540 614.600 ;
      RECT 927.500 1.400 927.780 614.600 ;
      RECT 929.740 1.400 930.020 614.600 ;
      RECT 931.980 1.400 932.260 614.600 ;
      RECT 934.220 1.400 934.500 614.600 ;
      RECT 936.460 1.400 936.740 614.600 ;
      RECT 938.700 1.400 938.980 614.600 ;
      RECT 940.940 1.400 941.220 614.600 ;
      RECT 943.180 1.400 943.460 614.600 ;
      RECT 945.420 1.400 945.700 614.600 ;
      RECT 947.660 1.400 947.940 614.600 ;
      RECT 949.900 1.400 950.180 614.600 ;
      RECT 952.140 1.400 952.420 614.600 ;
      RECT 954.380 1.400 954.660 614.600 ;
      RECT 956.620 1.400 956.900 614.600 ;
      RECT 958.860 1.400 959.140 614.600 ;
      RECT 961.100 1.400 961.380 614.600 ;
      RECT 963.340 1.400 963.620 614.600 ;
      RECT 965.580 1.400 965.860 614.600 ;
      RECT 967.820 1.400 968.100 614.600 ;
      RECT 970.060 1.400 970.340 614.600 ;
      RECT 972.300 1.400 972.580 614.600 ;
      RECT 974.540 1.400 974.820 614.600 ;
      RECT 976.780 1.400 977.060 614.600 ;
      RECT 979.020 1.400 979.300 614.600 ;
      RECT 981.260 1.400 981.540 614.600 ;
      RECT 983.500 1.400 983.780 614.600 ;
      RECT 985.740 1.400 986.020 614.600 ;
      RECT 987.980 1.400 988.260 614.600 ;
      RECT 990.220 1.400 990.500 614.600 ;
      RECT 992.460 1.400 992.740 614.600 ;
      RECT 994.700 1.400 994.980 614.600 ;
      RECT 996.940 1.400 997.220 614.600 ;
      RECT 999.180 1.400 999.460 614.600 ;
      RECT 1001.420 1.400 1001.700 614.600 ;
      RECT 1003.660 1.400 1003.940 614.600 ;
      RECT 1005.900 1.400 1006.180 614.600 ;
      RECT 1008.140 1.400 1008.420 614.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 1010.230 616.000 ;
    LAYER metal2 ;
    RECT 0 0 1010.230 616.000 ;
    LAYER metal3 ;
    RECT 0.070 0 1010.230 616.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 6.685 ;
    RECT 0 6.755 0.070 12.005 ;
    RECT 0 12.075 0.070 17.325 ;
    RECT 0 17.395 0.070 22.645 ;
    RECT 0 22.715 0.070 27.965 ;
    RECT 0 28.035 0.070 33.285 ;
    RECT 0 33.355 0.070 38.605 ;
    RECT 0 38.675 0.070 43.925 ;
    RECT 0 43.995 0.070 49.245 ;
    RECT 0 49.315 0.070 54.565 ;
    RECT 0 54.635 0.070 59.885 ;
    RECT 0 59.955 0.070 65.205 ;
    RECT 0 65.275 0.070 70.525 ;
    RECT 0 70.595 0.070 75.845 ;
    RECT 0 75.915 0.070 81.165 ;
    RECT 0 81.235 0.070 86.485 ;
    RECT 0 86.555 0.070 91.805 ;
    RECT 0 91.875 0.070 97.125 ;
    RECT 0 97.195 0.070 102.445 ;
    RECT 0 102.515 0.070 107.765 ;
    RECT 0 107.835 0.070 113.085 ;
    RECT 0 113.155 0.070 118.405 ;
    RECT 0 118.475 0.070 123.725 ;
    RECT 0 123.795 0.070 129.045 ;
    RECT 0 129.115 0.070 134.365 ;
    RECT 0 134.435 0.070 139.685 ;
    RECT 0 139.755 0.070 145.005 ;
    RECT 0 145.075 0.070 150.325 ;
    RECT 0 150.395 0.070 155.645 ;
    RECT 0 155.715 0.070 160.965 ;
    RECT 0 161.035 0.070 166.285 ;
    RECT 0 166.355 0.070 169.225 ;
    RECT 0 169.295 0.070 174.545 ;
    RECT 0 174.615 0.070 179.865 ;
    RECT 0 179.935 0.070 185.185 ;
    RECT 0 185.255 0.070 190.505 ;
    RECT 0 190.575 0.070 195.825 ;
    RECT 0 195.895 0.070 201.145 ;
    RECT 0 201.215 0.070 206.465 ;
    RECT 0 206.535 0.070 211.785 ;
    RECT 0 211.855 0.070 217.105 ;
    RECT 0 217.175 0.070 222.425 ;
    RECT 0 222.495 0.070 227.745 ;
    RECT 0 227.815 0.070 233.065 ;
    RECT 0 233.135 0.070 238.385 ;
    RECT 0 238.455 0.070 243.705 ;
    RECT 0 243.775 0.070 249.025 ;
    RECT 0 249.095 0.070 254.345 ;
    RECT 0 254.415 0.070 259.665 ;
    RECT 0 259.735 0.070 264.985 ;
    RECT 0 265.055 0.070 270.305 ;
    RECT 0 270.375 0.070 275.625 ;
    RECT 0 275.695 0.070 280.945 ;
    RECT 0 281.015 0.070 286.265 ;
    RECT 0 286.335 0.070 291.585 ;
    RECT 0 291.655 0.070 296.905 ;
    RECT 0 296.975 0.070 302.225 ;
    RECT 0 302.295 0.070 307.545 ;
    RECT 0 307.615 0.070 312.865 ;
    RECT 0 312.935 0.070 318.185 ;
    RECT 0 318.255 0.070 323.505 ;
    RECT 0 323.575 0.070 328.825 ;
    RECT 0 328.895 0.070 334.145 ;
    RECT 0 334.215 0.070 337.085 ;
    RECT 0 337.155 0.070 342.405 ;
    RECT 0 342.475 0.070 347.725 ;
    RECT 0 347.795 0.070 353.045 ;
    RECT 0 353.115 0.070 358.365 ;
    RECT 0 358.435 0.070 363.685 ;
    RECT 0 363.755 0.070 369.005 ;
    RECT 0 369.075 0.070 374.325 ;
    RECT 0 374.395 0.070 379.645 ;
    RECT 0 379.715 0.070 384.965 ;
    RECT 0 385.035 0.070 390.285 ;
    RECT 0 390.355 0.070 395.605 ;
    RECT 0 395.675 0.070 400.925 ;
    RECT 0 400.995 0.070 406.245 ;
    RECT 0 406.315 0.070 411.565 ;
    RECT 0 411.635 0.070 416.885 ;
    RECT 0 416.955 0.070 422.205 ;
    RECT 0 422.275 0.070 427.525 ;
    RECT 0 427.595 0.070 432.845 ;
    RECT 0 432.915 0.070 438.165 ;
    RECT 0 438.235 0.070 443.485 ;
    RECT 0 443.555 0.070 448.805 ;
    RECT 0 448.875 0.070 454.125 ;
    RECT 0 454.195 0.070 459.445 ;
    RECT 0 459.515 0.070 464.765 ;
    RECT 0 464.835 0.070 470.085 ;
    RECT 0 470.155 0.070 475.405 ;
    RECT 0 475.475 0.070 480.725 ;
    RECT 0 480.795 0.070 486.045 ;
    RECT 0 486.115 0.070 491.365 ;
    RECT 0 491.435 0.070 496.685 ;
    RECT 0 496.755 0.070 502.005 ;
    RECT 0 502.075 0.070 504.945 ;
    RECT 0 505.015 0.070 510.265 ;
    RECT 0 510.335 0.070 515.585 ;
    RECT 0 515.655 0.070 520.905 ;
    RECT 0 520.975 0.070 526.225 ;
    RECT 0 526.295 0.070 531.545 ;
    RECT 0 531.615 0.070 536.865 ;
    RECT 0 536.935 0.070 542.185 ;
    RECT 0 542.255 0.070 547.505 ;
    RECT 0 547.575 0.070 552.825 ;
    RECT 0 552.895 0.070 558.145 ;
    RECT 0 558.215 0.070 563.465 ;
    RECT 0 563.535 0.070 568.785 ;
    RECT 0 568.855 0.070 574.105 ;
    RECT 0 574.175 0.070 577.045 ;
    RECT 0 577.115 0.070 582.365 ;
    RECT 0 582.435 0.070 587.685 ;
    RECT 0 587.755 0.070 616.000 ;
    LAYER metal4 ;
    RECT 0 0 1010.230 1.400 ;
    RECT 0 614.600 1010.230 616.000 ;
    RECT 0.000 1.400 1.260 614.600 ;
    RECT 1.540 1.400 2.380 614.600 ;
    RECT 2.660 1.400 3.500 614.600 ;
    RECT 3.780 1.400 4.620 614.600 ;
    RECT 4.900 1.400 5.740 614.600 ;
    RECT 6.020 1.400 6.860 614.600 ;
    RECT 7.140 1.400 7.980 614.600 ;
    RECT 8.260 1.400 9.100 614.600 ;
    RECT 9.380 1.400 10.220 614.600 ;
    RECT 10.500 1.400 11.340 614.600 ;
    RECT 11.620 1.400 12.460 614.600 ;
    RECT 12.740 1.400 13.580 614.600 ;
    RECT 13.860 1.400 14.700 614.600 ;
    RECT 14.980 1.400 15.820 614.600 ;
    RECT 16.100 1.400 16.940 614.600 ;
    RECT 17.220 1.400 18.060 614.600 ;
    RECT 18.340 1.400 19.180 614.600 ;
    RECT 19.460 1.400 20.300 614.600 ;
    RECT 20.580 1.400 21.420 614.600 ;
    RECT 21.700 1.400 22.540 614.600 ;
    RECT 22.820 1.400 23.660 614.600 ;
    RECT 23.940 1.400 24.780 614.600 ;
    RECT 25.060 1.400 25.900 614.600 ;
    RECT 26.180 1.400 27.020 614.600 ;
    RECT 27.300 1.400 28.140 614.600 ;
    RECT 28.420 1.400 29.260 614.600 ;
    RECT 29.540 1.400 30.380 614.600 ;
    RECT 30.660 1.400 31.500 614.600 ;
    RECT 31.780 1.400 32.620 614.600 ;
    RECT 32.900 1.400 33.740 614.600 ;
    RECT 34.020 1.400 34.860 614.600 ;
    RECT 35.140 1.400 35.980 614.600 ;
    RECT 36.260 1.400 37.100 614.600 ;
    RECT 37.380 1.400 38.220 614.600 ;
    RECT 38.500 1.400 39.340 614.600 ;
    RECT 39.620 1.400 40.460 614.600 ;
    RECT 40.740 1.400 41.580 614.600 ;
    RECT 41.860 1.400 42.700 614.600 ;
    RECT 42.980 1.400 43.820 614.600 ;
    RECT 44.100 1.400 44.940 614.600 ;
    RECT 45.220 1.400 46.060 614.600 ;
    RECT 46.340 1.400 47.180 614.600 ;
    RECT 47.460 1.400 48.300 614.600 ;
    RECT 48.580 1.400 49.420 614.600 ;
    RECT 49.700 1.400 50.540 614.600 ;
    RECT 50.820 1.400 51.660 614.600 ;
    RECT 51.940 1.400 52.780 614.600 ;
    RECT 53.060 1.400 53.900 614.600 ;
    RECT 54.180 1.400 55.020 614.600 ;
    RECT 55.300 1.400 56.140 614.600 ;
    RECT 56.420 1.400 57.260 614.600 ;
    RECT 57.540 1.400 58.380 614.600 ;
    RECT 58.660 1.400 59.500 614.600 ;
    RECT 59.780 1.400 60.620 614.600 ;
    RECT 60.900 1.400 61.740 614.600 ;
    RECT 62.020 1.400 62.860 614.600 ;
    RECT 63.140 1.400 63.980 614.600 ;
    RECT 64.260 1.400 65.100 614.600 ;
    RECT 65.380 1.400 66.220 614.600 ;
    RECT 66.500 1.400 67.340 614.600 ;
    RECT 67.620 1.400 68.460 614.600 ;
    RECT 68.740 1.400 69.580 614.600 ;
    RECT 69.860 1.400 70.700 614.600 ;
    RECT 70.980 1.400 71.820 614.600 ;
    RECT 72.100 1.400 72.940 614.600 ;
    RECT 73.220 1.400 74.060 614.600 ;
    RECT 74.340 1.400 75.180 614.600 ;
    RECT 75.460 1.400 76.300 614.600 ;
    RECT 76.580 1.400 77.420 614.600 ;
    RECT 77.700 1.400 78.540 614.600 ;
    RECT 78.820 1.400 79.660 614.600 ;
    RECT 79.940 1.400 80.780 614.600 ;
    RECT 81.060 1.400 81.900 614.600 ;
    RECT 82.180 1.400 83.020 614.600 ;
    RECT 83.300 1.400 84.140 614.600 ;
    RECT 84.420 1.400 85.260 614.600 ;
    RECT 85.540 1.400 86.380 614.600 ;
    RECT 86.660 1.400 87.500 614.600 ;
    RECT 87.780 1.400 88.620 614.600 ;
    RECT 88.900 1.400 89.740 614.600 ;
    RECT 90.020 1.400 90.860 614.600 ;
    RECT 91.140 1.400 91.980 614.600 ;
    RECT 92.260 1.400 93.100 614.600 ;
    RECT 93.380 1.400 94.220 614.600 ;
    RECT 94.500 1.400 95.340 614.600 ;
    RECT 95.620 1.400 96.460 614.600 ;
    RECT 96.740 1.400 97.580 614.600 ;
    RECT 97.860 1.400 98.700 614.600 ;
    RECT 98.980 1.400 99.820 614.600 ;
    RECT 100.100 1.400 100.940 614.600 ;
    RECT 101.220 1.400 102.060 614.600 ;
    RECT 102.340 1.400 103.180 614.600 ;
    RECT 103.460 1.400 104.300 614.600 ;
    RECT 104.580 1.400 105.420 614.600 ;
    RECT 105.700 1.400 106.540 614.600 ;
    RECT 106.820 1.400 107.660 614.600 ;
    RECT 107.940 1.400 108.780 614.600 ;
    RECT 109.060 1.400 109.900 614.600 ;
    RECT 110.180 1.400 111.020 614.600 ;
    RECT 111.300 1.400 112.140 614.600 ;
    RECT 112.420 1.400 113.260 614.600 ;
    RECT 113.540 1.400 114.380 614.600 ;
    RECT 114.660 1.400 115.500 614.600 ;
    RECT 115.780 1.400 116.620 614.600 ;
    RECT 116.900 1.400 117.740 614.600 ;
    RECT 118.020 1.400 118.860 614.600 ;
    RECT 119.140 1.400 119.980 614.600 ;
    RECT 120.260 1.400 121.100 614.600 ;
    RECT 121.380 1.400 122.220 614.600 ;
    RECT 122.500 1.400 123.340 614.600 ;
    RECT 123.620 1.400 124.460 614.600 ;
    RECT 124.740 1.400 125.580 614.600 ;
    RECT 125.860 1.400 126.700 614.600 ;
    RECT 126.980 1.400 127.820 614.600 ;
    RECT 128.100 1.400 128.940 614.600 ;
    RECT 129.220 1.400 130.060 614.600 ;
    RECT 130.340 1.400 131.180 614.600 ;
    RECT 131.460 1.400 132.300 614.600 ;
    RECT 132.580 1.400 133.420 614.600 ;
    RECT 133.700 1.400 134.540 614.600 ;
    RECT 134.820 1.400 135.660 614.600 ;
    RECT 135.940 1.400 136.780 614.600 ;
    RECT 137.060 1.400 137.900 614.600 ;
    RECT 138.180 1.400 139.020 614.600 ;
    RECT 139.300 1.400 140.140 614.600 ;
    RECT 140.420 1.400 141.260 614.600 ;
    RECT 141.540 1.400 142.380 614.600 ;
    RECT 142.660 1.400 143.500 614.600 ;
    RECT 143.780 1.400 144.620 614.600 ;
    RECT 144.900 1.400 145.740 614.600 ;
    RECT 146.020 1.400 146.860 614.600 ;
    RECT 147.140 1.400 147.980 614.600 ;
    RECT 148.260 1.400 149.100 614.600 ;
    RECT 149.380 1.400 150.220 614.600 ;
    RECT 150.500 1.400 151.340 614.600 ;
    RECT 151.620 1.400 152.460 614.600 ;
    RECT 152.740 1.400 153.580 614.600 ;
    RECT 153.860 1.400 154.700 614.600 ;
    RECT 154.980 1.400 155.820 614.600 ;
    RECT 156.100 1.400 156.940 614.600 ;
    RECT 157.220 1.400 158.060 614.600 ;
    RECT 158.340 1.400 159.180 614.600 ;
    RECT 159.460 1.400 160.300 614.600 ;
    RECT 160.580 1.400 161.420 614.600 ;
    RECT 161.700 1.400 162.540 614.600 ;
    RECT 162.820 1.400 163.660 614.600 ;
    RECT 163.940 1.400 164.780 614.600 ;
    RECT 165.060 1.400 165.900 614.600 ;
    RECT 166.180 1.400 167.020 614.600 ;
    RECT 167.300 1.400 168.140 614.600 ;
    RECT 168.420 1.400 169.260 614.600 ;
    RECT 169.540 1.400 170.380 614.600 ;
    RECT 170.660 1.400 171.500 614.600 ;
    RECT 171.780 1.400 172.620 614.600 ;
    RECT 172.900 1.400 173.740 614.600 ;
    RECT 174.020 1.400 174.860 614.600 ;
    RECT 175.140 1.400 175.980 614.600 ;
    RECT 176.260 1.400 177.100 614.600 ;
    RECT 177.380 1.400 178.220 614.600 ;
    RECT 178.500 1.400 179.340 614.600 ;
    RECT 179.620 1.400 180.460 614.600 ;
    RECT 180.740 1.400 181.580 614.600 ;
    RECT 181.860 1.400 182.700 614.600 ;
    RECT 182.980 1.400 183.820 614.600 ;
    RECT 184.100 1.400 184.940 614.600 ;
    RECT 185.220 1.400 186.060 614.600 ;
    RECT 186.340 1.400 187.180 614.600 ;
    RECT 187.460 1.400 188.300 614.600 ;
    RECT 188.580 1.400 189.420 614.600 ;
    RECT 189.700 1.400 190.540 614.600 ;
    RECT 190.820 1.400 191.660 614.600 ;
    RECT 191.940 1.400 192.780 614.600 ;
    RECT 193.060 1.400 193.900 614.600 ;
    RECT 194.180 1.400 195.020 614.600 ;
    RECT 195.300 1.400 196.140 614.600 ;
    RECT 196.420 1.400 197.260 614.600 ;
    RECT 197.540 1.400 198.380 614.600 ;
    RECT 198.660 1.400 199.500 614.600 ;
    RECT 199.780 1.400 200.620 614.600 ;
    RECT 200.900 1.400 201.740 614.600 ;
    RECT 202.020 1.400 202.860 614.600 ;
    RECT 203.140 1.400 203.980 614.600 ;
    RECT 204.260 1.400 205.100 614.600 ;
    RECT 205.380 1.400 206.220 614.600 ;
    RECT 206.500 1.400 207.340 614.600 ;
    RECT 207.620 1.400 208.460 614.600 ;
    RECT 208.740 1.400 209.580 614.600 ;
    RECT 209.860 1.400 210.700 614.600 ;
    RECT 210.980 1.400 211.820 614.600 ;
    RECT 212.100 1.400 212.940 614.600 ;
    RECT 213.220 1.400 214.060 614.600 ;
    RECT 214.340 1.400 215.180 614.600 ;
    RECT 215.460 1.400 216.300 614.600 ;
    RECT 216.580 1.400 217.420 614.600 ;
    RECT 217.700 1.400 218.540 614.600 ;
    RECT 218.820 1.400 219.660 614.600 ;
    RECT 219.940 1.400 220.780 614.600 ;
    RECT 221.060 1.400 221.900 614.600 ;
    RECT 222.180 1.400 223.020 614.600 ;
    RECT 223.300 1.400 224.140 614.600 ;
    RECT 224.420 1.400 225.260 614.600 ;
    RECT 225.540 1.400 226.380 614.600 ;
    RECT 226.660 1.400 227.500 614.600 ;
    RECT 227.780 1.400 228.620 614.600 ;
    RECT 228.900 1.400 229.740 614.600 ;
    RECT 230.020 1.400 230.860 614.600 ;
    RECT 231.140 1.400 231.980 614.600 ;
    RECT 232.260 1.400 233.100 614.600 ;
    RECT 233.380 1.400 234.220 614.600 ;
    RECT 234.500 1.400 235.340 614.600 ;
    RECT 235.620 1.400 236.460 614.600 ;
    RECT 236.740 1.400 237.580 614.600 ;
    RECT 237.860 1.400 238.700 614.600 ;
    RECT 238.980 1.400 239.820 614.600 ;
    RECT 240.100 1.400 240.940 614.600 ;
    RECT 241.220 1.400 242.060 614.600 ;
    RECT 242.340 1.400 243.180 614.600 ;
    RECT 243.460 1.400 244.300 614.600 ;
    RECT 244.580 1.400 245.420 614.600 ;
    RECT 245.700 1.400 246.540 614.600 ;
    RECT 246.820 1.400 247.660 614.600 ;
    RECT 247.940 1.400 248.780 614.600 ;
    RECT 249.060 1.400 249.900 614.600 ;
    RECT 250.180 1.400 251.020 614.600 ;
    RECT 251.300 1.400 252.140 614.600 ;
    RECT 252.420 1.400 253.260 614.600 ;
    RECT 253.540 1.400 254.380 614.600 ;
    RECT 254.660 1.400 255.500 614.600 ;
    RECT 255.780 1.400 256.620 614.600 ;
    RECT 256.900 1.400 257.740 614.600 ;
    RECT 258.020 1.400 258.860 614.600 ;
    RECT 259.140 1.400 259.980 614.600 ;
    RECT 260.260 1.400 261.100 614.600 ;
    RECT 261.380 1.400 262.220 614.600 ;
    RECT 262.500 1.400 263.340 614.600 ;
    RECT 263.620 1.400 264.460 614.600 ;
    RECT 264.740 1.400 265.580 614.600 ;
    RECT 265.860 1.400 266.700 614.600 ;
    RECT 266.980 1.400 267.820 614.600 ;
    RECT 268.100 1.400 268.940 614.600 ;
    RECT 269.220 1.400 270.060 614.600 ;
    RECT 270.340 1.400 271.180 614.600 ;
    RECT 271.460 1.400 272.300 614.600 ;
    RECT 272.580 1.400 273.420 614.600 ;
    RECT 273.700 1.400 274.540 614.600 ;
    RECT 274.820 1.400 275.660 614.600 ;
    RECT 275.940 1.400 276.780 614.600 ;
    RECT 277.060 1.400 277.900 614.600 ;
    RECT 278.180 1.400 279.020 614.600 ;
    RECT 279.300 1.400 280.140 614.600 ;
    RECT 280.420 1.400 281.260 614.600 ;
    RECT 281.540 1.400 282.380 614.600 ;
    RECT 282.660 1.400 283.500 614.600 ;
    RECT 283.780 1.400 284.620 614.600 ;
    RECT 284.900 1.400 285.740 614.600 ;
    RECT 286.020 1.400 286.860 614.600 ;
    RECT 287.140 1.400 287.980 614.600 ;
    RECT 288.260 1.400 289.100 614.600 ;
    RECT 289.380 1.400 290.220 614.600 ;
    RECT 290.500 1.400 291.340 614.600 ;
    RECT 291.620 1.400 292.460 614.600 ;
    RECT 292.740 1.400 293.580 614.600 ;
    RECT 293.860 1.400 294.700 614.600 ;
    RECT 294.980 1.400 295.820 614.600 ;
    RECT 296.100 1.400 296.940 614.600 ;
    RECT 297.220 1.400 298.060 614.600 ;
    RECT 298.340 1.400 299.180 614.600 ;
    RECT 299.460 1.400 300.300 614.600 ;
    RECT 300.580 1.400 301.420 614.600 ;
    RECT 301.700 1.400 302.540 614.600 ;
    RECT 302.820 1.400 303.660 614.600 ;
    RECT 303.940 1.400 304.780 614.600 ;
    RECT 305.060 1.400 305.900 614.600 ;
    RECT 306.180 1.400 307.020 614.600 ;
    RECT 307.300 1.400 308.140 614.600 ;
    RECT 308.420 1.400 309.260 614.600 ;
    RECT 309.540 1.400 310.380 614.600 ;
    RECT 310.660 1.400 311.500 614.600 ;
    RECT 311.780 1.400 312.620 614.600 ;
    RECT 312.900 1.400 313.740 614.600 ;
    RECT 314.020 1.400 314.860 614.600 ;
    RECT 315.140 1.400 315.980 614.600 ;
    RECT 316.260 1.400 317.100 614.600 ;
    RECT 317.380 1.400 318.220 614.600 ;
    RECT 318.500 1.400 319.340 614.600 ;
    RECT 319.620 1.400 320.460 614.600 ;
    RECT 320.740 1.400 321.580 614.600 ;
    RECT 321.860 1.400 322.700 614.600 ;
    RECT 322.980 1.400 323.820 614.600 ;
    RECT 324.100 1.400 324.940 614.600 ;
    RECT 325.220 1.400 326.060 614.600 ;
    RECT 326.340 1.400 327.180 614.600 ;
    RECT 327.460 1.400 328.300 614.600 ;
    RECT 328.580 1.400 329.420 614.600 ;
    RECT 329.700 1.400 330.540 614.600 ;
    RECT 330.820 1.400 331.660 614.600 ;
    RECT 331.940 1.400 332.780 614.600 ;
    RECT 333.060 1.400 333.900 614.600 ;
    RECT 334.180 1.400 335.020 614.600 ;
    RECT 335.300 1.400 336.140 614.600 ;
    RECT 336.420 1.400 337.260 614.600 ;
    RECT 337.540 1.400 338.380 614.600 ;
    RECT 338.660 1.400 339.500 614.600 ;
    RECT 339.780 1.400 340.620 614.600 ;
    RECT 340.900 1.400 341.740 614.600 ;
    RECT 342.020 1.400 342.860 614.600 ;
    RECT 343.140 1.400 343.980 614.600 ;
    RECT 344.260 1.400 345.100 614.600 ;
    RECT 345.380 1.400 346.220 614.600 ;
    RECT 346.500 1.400 347.340 614.600 ;
    RECT 347.620 1.400 348.460 614.600 ;
    RECT 348.740 1.400 349.580 614.600 ;
    RECT 349.860 1.400 350.700 614.600 ;
    RECT 350.980 1.400 351.820 614.600 ;
    RECT 352.100 1.400 352.940 614.600 ;
    RECT 353.220 1.400 354.060 614.600 ;
    RECT 354.340 1.400 355.180 614.600 ;
    RECT 355.460 1.400 356.300 614.600 ;
    RECT 356.580 1.400 357.420 614.600 ;
    RECT 357.700 1.400 358.540 614.600 ;
    RECT 358.820 1.400 359.660 614.600 ;
    RECT 359.940 1.400 360.780 614.600 ;
    RECT 361.060 1.400 361.900 614.600 ;
    RECT 362.180 1.400 363.020 614.600 ;
    RECT 363.300 1.400 364.140 614.600 ;
    RECT 364.420 1.400 365.260 614.600 ;
    RECT 365.540 1.400 366.380 614.600 ;
    RECT 366.660 1.400 367.500 614.600 ;
    RECT 367.780 1.400 368.620 614.600 ;
    RECT 368.900 1.400 369.740 614.600 ;
    RECT 370.020 1.400 370.860 614.600 ;
    RECT 371.140 1.400 371.980 614.600 ;
    RECT 372.260 1.400 373.100 614.600 ;
    RECT 373.380 1.400 374.220 614.600 ;
    RECT 374.500 1.400 375.340 614.600 ;
    RECT 375.620 1.400 376.460 614.600 ;
    RECT 376.740 1.400 377.580 614.600 ;
    RECT 377.860 1.400 378.700 614.600 ;
    RECT 378.980 1.400 379.820 614.600 ;
    RECT 380.100 1.400 380.940 614.600 ;
    RECT 381.220 1.400 382.060 614.600 ;
    RECT 382.340 1.400 383.180 614.600 ;
    RECT 383.460 1.400 384.300 614.600 ;
    RECT 384.580 1.400 385.420 614.600 ;
    RECT 385.700 1.400 386.540 614.600 ;
    RECT 386.820 1.400 387.660 614.600 ;
    RECT 387.940 1.400 388.780 614.600 ;
    RECT 389.060 1.400 389.900 614.600 ;
    RECT 390.180 1.400 391.020 614.600 ;
    RECT 391.300 1.400 392.140 614.600 ;
    RECT 392.420 1.400 393.260 614.600 ;
    RECT 393.540 1.400 394.380 614.600 ;
    RECT 394.660 1.400 395.500 614.600 ;
    RECT 395.780 1.400 396.620 614.600 ;
    RECT 396.900 1.400 397.740 614.600 ;
    RECT 398.020 1.400 398.860 614.600 ;
    RECT 399.140 1.400 399.980 614.600 ;
    RECT 400.260 1.400 401.100 614.600 ;
    RECT 401.380 1.400 402.220 614.600 ;
    RECT 402.500 1.400 403.340 614.600 ;
    RECT 403.620 1.400 404.460 614.600 ;
    RECT 404.740 1.400 405.580 614.600 ;
    RECT 405.860 1.400 406.700 614.600 ;
    RECT 406.980 1.400 407.820 614.600 ;
    RECT 408.100 1.400 408.940 614.600 ;
    RECT 409.220 1.400 410.060 614.600 ;
    RECT 410.340 1.400 411.180 614.600 ;
    RECT 411.460 1.400 412.300 614.600 ;
    RECT 412.580 1.400 413.420 614.600 ;
    RECT 413.700 1.400 414.540 614.600 ;
    RECT 414.820 1.400 415.660 614.600 ;
    RECT 415.940 1.400 416.780 614.600 ;
    RECT 417.060 1.400 417.900 614.600 ;
    RECT 418.180 1.400 419.020 614.600 ;
    RECT 419.300 1.400 420.140 614.600 ;
    RECT 420.420 1.400 421.260 614.600 ;
    RECT 421.540 1.400 422.380 614.600 ;
    RECT 422.660 1.400 423.500 614.600 ;
    RECT 423.780 1.400 424.620 614.600 ;
    RECT 424.900 1.400 425.740 614.600 ;
    RECT 426.020 1.400 426.860 614.600 ;
    RECT 427.140 1.400 427.980 614.600 ;
    RECT 428.260 1.400 429.100 614.600 ;
    RECT 429.380 1.400 430.220 614.600 ;
    RECT 430.500 1.400 431.340 614.600 ;
    RECT 431.620 1.400 432.460 614.600 ;
    RECT 432.740 1.400 433.580 614.600 ;
    RECT 433.860 1.400 434.700 614.600 ;
    RECT 434.980 1.400 435.820 614.600 ;
    RECT 436.100 1.400 436.940 614.600 ;
    RECT 437.220 1.400 438.060 614.600 ;
    RECT 438.340 1.400 439.180 614.600 ;
    RECT 439.460 1.400 440.300 614.600 ;
    RECT 440.580 1.400 441.420 614.600 ;
    RECT 441.700 1.400 442.540 614.600 ;
    RECT 442.820 1.400 443.660 614.600 ;
    RECT 443.940 1.400 444.780 614.600 ;
    RECT 445.060 1.400 445.900 614.600 ;
    RECT 446.180 1.400 447.020 614.600 ;
    RECT 447.300 1.400 448.140 614.600 ;
    RECT 448.420 1.400 449.260 614.600 ;
    RECT 449.540 1.400 450.380 614.600 ;
    RECT 450.660 1.400 451.500 614.600 ;
    RECT 451.780 1.400 452.620 614.600 ;
    RECT 452.900 1.400 453.740 614.600 ;
    RECT 454.020 1.400 454.860 614.600 ;
    RECT 455.140 1.400 455.980 614.600 ;
    RECT 456.260 1.400 457.100 614.600 ;
    RECT 457.380 1.400 458.220 614.600 ;
    RECT 458.500 1.400 459.340 614.600 ;
    RECT 459.620 1.400 460.460 614.600 ;
    RECT 460.740 1.400 461.580 614.600 ;
    RECT 461.860 1.400 462.700 614.600 ;
    RECT 462.980 1.400 463.820 614.600 ;
    RECT 464.100 1.400 464.940 614.600 ;
    RECT 465.220 1.400 466.060 614.600 ;
    RECT 466.340 1.400 467.180 614.600 ;
    RECT 467.460 1.400 468.300 614.600 ;
    RECT 468.580 1.400 469.420 614.600 ;
    RECT 469.700 1.400 470.540 614.600 ;
    RECT 470.820 1.400 471.660 614.600 ;
    RECT 471.940 1.400 472.780 614.600 ;
    RECT 473.060 1.400 473.900 614.600 ;
    RECT 474.180 1.400 475.020 614.600 ;
    RECT 475.300 1.400 476.140 614.600 ;
    RECT 476.420 1.400 477.260 614.600 ;
    RECT 477.540 1.400 478.380 614.600 ;
    RECT 478.660 1.400 479.500 614.600 ;
    RECT 479.780 1.400 480.620 614.600 ;
    RECT 480.900 1.400 481.740 614.600 ;
    RECT 482.020 1.400 482.860 614.600 ;
    RECT 483.140 1.400 483.980 614.600 ;
    RECT 484.260 1.400 485.100 614.600 ;
    RECT 485.380 1.400 486.220 614.600 ;
    RECT 486.500 1.400 487.340 614.600 ;
    RECT 487.620 1.400 488.460 614.600 ;
    RECT 488.740 1.400 489.580 614.600 ;
    RECT 489.860 1.400 490.700 614.600 ;
    RECT 490.980 1.400 491.820 614.600 ;
    RECT 492.100 1.400 492.940 614.600 ;
    RECT 493.220 1.400 494.060 614.600 ;
    RECT 494.340 1.400 495.180 614.600 ;
    RECT 495.460 1.400 496.300 614.600 ;
    RECT 496.580 1.400 497.420 614.600 ;
    RECT 497.700 1.400 498.540 614.600 ;
    RECT 498.820 1.400 499.660 614.600 ;
    RECT 499.940 1.400 500.780 614.600 ;
    RECT 501.060 1.400 501.900 614.600 ;
    RECT 502.180 1.400 503.020 614.600 ;
    RECT 503.300 1.400 504.140 614.600 ;
    RECT 504.420 1.400 505.260 614.600 ;
    RECT 505.540 1.400 506.380 614.600 ;
    RECT 506.660 1.400 507.500 614.600 ;
    RECT 507.780 1.400 508.620 614.600 ;
    RECT 508.900 1.400 509.740 614.600 ;
    RECT 510.020 1.400 510.860 614.600 ;
    RECT 511.140 1.400 511.980 614.600 ;
    RECT 512.260 1.400 513.100 614.600 ;
    RECT 513.380 1.400 514.220 614.600 ;
    RECT 514.500 1.400 515.340 614.600 ;
    RECT 515.620 1.400 516.460 614.600 ;
    RECT 516.740 1.400 517.580 614.600 ;
    RECT 517.860 1.400 518.700 614.600 ;
    RECT 518.980 1.400 519.820 614.600 ;
    RECT 520.100 1.400 520.940 614.600 ;
    RECT 521.220 1.400 522.060 614.600 ;
    RECT 522.340 1.400 523.180 614.600 ;
    RECT 523.460 1.400 524.300 614.600 ;
    RECT 524.580 1.400 525.420 614.600 ;
    RECT 525.700 1.400 526.540 614.600 ;
    RECT 526.820 1.400 527.660 614.600 ;
    RECT 527.940 1.400 528.780 614.600 ;
    RECT 529.060 1.400 529.900 614.600 ;
    RECT 530.180 1.400 531.020 614.600 ;
    RECT 531.300 1.400 532.140 614.600 ;
    RECT 532.420 1.400 533.260 614.600 ;
    RECT 533.540 1.400 534.380 614.600 ;
    RECT 534.660 1.400 535.500 614.600 ;
    RECT 535.780 1.400 536.620 614.600 ;
    RECT 536.900 1.400 537.740 614.600 ;
    RECT 538.020 1.400 538.860 614.600 ;
    RECT 539.140 1.400 539.980 614.600 ;
    RECT 540.260 1.400 541.100 614.600 ;
    RECT 541.380 1.400 542.220 614.600 ;
    RECT 542.500 1.400 543.340 614.600 ;
    RECT 543.620 1.400 544.460 614.600 ;
    RECT 544.740 1.400 545.580 614.600 ;
    RECT 545.860 1.400 546.700 614.600 ;
    RECT 546.980 1.400 547.820 614.600 ;
    RECT 548.100 1.400 548.940 614.600 ;
    RECT 549.220 1.400 550.060 614.600 ;
    RECT 550.340 1.400 551.180 614.600 ;
    RECT 551.460 1.400 552.300 614.600 ;
    RECT 552.580 1.400 553.420 614.600 ;
    RECT 553.700 1.400 554.540 614.600 ;
    RECT 554.820 1.400 555.660 614.600 ;
    RECT 555.940 1.400 556.780 614.600 ;
    RECT 557.060 1.400 557.900 614.600 ;
    RECT 558.180 1.400 559.020 614.600 ;
    RECT 559.300 1.400 560.140 614.600 ;
    RECT 560.420 1.400 561.260 614.600 ;
    RECT 561.540 1.400 562.380 614.600 ;
    RECT 562.660 1.400 563.500 614.600 ;
    RECT 563.780 1.400 564.620 614.600 ;
    RECT 564.900 1.400 565.740 614.600 ;
    RECT 566.020 1.400 566.860 614.600 ;
    RECT 567.140 1.400 567.980 614.600 ;
    RECT 568.260 1.400 569.100 614.600 ;
    RECT 569.380 1.400 570.220 614.600 ;
    RECT 570.500 1.400 571.340 614.600 ;
    RECT 571.620 1.400 572.460 614.600 ;
    RECT 572.740 1.400 573.580 614.600 ;
    RECT 573.860 1.400 574.700 614.600 ;
    RECT 574.980 1.400 575.820 614.600 ;
    RECT 576.100 1.400 576.940 614.600 ;
    RECT 577.220 1.400 578.060 614.600 ;
    RECT 578.340 1.400 579.180 614.600 ;
    RECT 579.460 1.400 580.300 614.600 ;
    RECT 580.580 1.400 581.420 614.600 ;
    RECT 581.700 1.400 582.540 614.600 ;
    RECT 582.820 1.400 583.660 614.600 ;
    RECT 583.940 1.400 584.780 614.600 ;
    RECT 585.060 1.400 585.900 614.600 ;
    RECT 586.180 1.400 587.020 614.600 ;
    RECT 587.300 1.400 588.140 614.600 ;
    RECT 588.420 1.400 589.260 614.600 ;
    RECT 589.540 1.400 590.380 614.600 ;
    RECT 590.660 1.400 591.500 614.600 ;
    RECT 591.780 1.400 592.620 614.600 ;
    RECT 592.900 1.400 593.740 614.600 ;
    RECT 594.020 1.400 594.860 614.600 ;
    RECT 595.140 1.400 595.980 614.600 ;
    RECT 596.260 1.400 597.100 614.600 ;
    RECT 597.380 1.400 598.220 614.600 ;
    RECT 598.500 1.400 599.340 614.600 ;
    RECT 599.620 1.400 600.460 614.600 ;
    RECT 600.740 1.400 601.580 614.600 ;
    RECT 601.860 1.400 602.700 614.600 ;
    RECT 602.980 1.400 603.820 614.600 ;
    RECT 604.100 1.400 604.940 614.600 ;
    RECT 605.220 1.400 606.060 614.600 ;
    RECT 606.340 1.400 607.180 614.600 ;
    RECT 607.460 1.400 608.300 614.600 ;
    RECT 608.580 1.400 609.420 614.600 ;
    RECT 609.700 1.400 610.540 614.600 ;
    RECT 610.820 1.400 611.660 614.600 ;
    RECT 611.940 1.400 612.780 614.600 ;
    RECT 613.060 1.400 613.900 614.600 ;
    RECT 614.180 1.400 615.020 614.600 ;
    RECT 615.300 1.400 616.140 614.600 ;
    RECT 616.420 1.400 617.260 614.600 ;
    RECT 617.540 1.400 618.380 614.600 ;
    RECT 618.660 1.400 619.500 614.600 ;
    RECT 619.780 1.400 620.620 614.600 ;
    RECT 620.900 1.400 621.740 614.600 ;
    RECT 622.020 1.400 622.860 614.600 ;
    RECT 623.140 1.400 623.980 614.600 ;
    RECT 624.260 1.400 625.100 614.600 ;
    RECT 625.380 1.400 626.220 614.600 ;
    RECT 626.500 1.400 627.340 614.600 ;
    RECT 627.620 1.400 628.460 614.600 ;
    RECT 628.740 1.400 629.580 614.600 ;
    RECT 629.860 1.400 630.700 614.600 ;
    RECT 630.980 1.400 631.820 614.600 ;
    RECT 632.100 1.400 632.940 614.600 ;
    RECT 633.220 1.400 634.060 614.600 ;
    RECT 634.340 1.400 635.180 614.600 ;
    RECT 635.460 1.400 636.300 614.600 ;
    RECT 636.580 1.400 637.420 614.600 ;
    RECT 637.700 1.400 638.540 614.600 ;
    RECT 638.820 1.400 639.660 614.600 ;
    RECT 639.940 1.400 640.780 614.600 ;
    RECT 641.060 1.400 641.900 614.600 ;
    RECT 642.180 1.400 643.020 614.600 ;
    RECT 643.300 1.400 644.140 614.600 ;
    RECT 644.420 1.400 645.260 614.600 ;
    RECT 645.540 1.400 646.380 614.600 ;
    RECT 646.660 1.400 647.500 614.600 ;
    RECT 647.780 1.400 648.620 614.600 ;
    RECT 648.900 1.400 649.740 614.600 ;
    RECT 650.020 1.400 650.860 614.600 ;
    RECT 651.140 1.400 651.980 614.600 ;
    RECT 652.260 1.400 653.100 614.600 ;
    RECT 653.380 1.400 654.220 614.600 ;
    RECT 654.500 1.400 655.340 614.600 ;
    RECT 655.620 1.400 656.460 614.600 ;
    RECT 656.740 1.400 657.580 614.600 ;
    RECT 657.860 1.400 658.700 614.600 ;
    RECT 658.980 1.400 659.820 614.600 ;
    RECT 660.100 1.400 660.940 614.600 ;
    RECT 661.220 1.400 662.060 614.600 ;
    RECT 662.340 1.400 663.180 614.600 ;
    RECT 663.460 1.400 664.300 614.600 ;
    RECT 664.580 1.400 665.420 614.600 ;
    RECT 665.700 1.400 666.540 614.600 ;
    RECT 666.820 1.400 667.660 614.600 ;
    RECT 667.940 1.400 668.780 614.600 ;
    RECT 669.060 1.400 669.900 614.600 ;
    RECT 670.180 1.400 671.020 614.600 ;
    RECT 671.300 1.400 672.140 614.600 ;
    RECT 672.420 1.400 673.260 614.600 ;
    RECT 673.540 1.400 674.380 614.600 ;
    RECT 674.660 1.400 675.500 614.600 ;
    RECT 675.780 1.400 676.620 614.600 ;
    RECT 676.900 1.400 677.740 614.600 ;
    RECT 678.020 1.400 678.860 614.600 ;
    RECT 679.140 1.400 679.980 614.600 ;
    RECT 680.260 1.400 681.100 614.600 ;
    RECT 681.380 1.400 682.220 614.600 ;
    RECT 682.500 1.400 683.340 614.600 ;
    RECT 683.620 1.400 684.460 614.600 ;
    RECT 684.740 1.400 685.580 614.600 ;
    RECT 685.860 1.400 686.700 614.600 ;
    RECT 686.980 1.400 687.820 614.600 ;
    RECT 688.100 1.400 688.940 614.600 ;
    RECT 689.220 1.400 690.060 614.600 ;
    RECT 690.340 1.400 691.180 614.600 ;
    RECT 691.460 1.400 692.300 614.600 ;
    RECT 692.580 1.400 693.420 614.600 ;
    RECT 693.700 1.400 694.540 614.600 ;
    RECT 694.820 1.400 695.660 614.600 ;
    RECT 695.940 1.400 696.780 614.600 ;
    RECT 697.060 1.400 697.900 614.600 ;
    RECT 698.180 1.400 699.020 614.600 ;
    RECT 699.300 1.400 700.140 614.600 ;
    RECT 700.420 1.400 701.260 614.600 ;
    RECT 701.540 1.400 702.380 614.600 ;
    RECT 702.660 1.400 703.500 614.600 ;
    RECT 703.780 1.400 704.620 614.600 ;
    RECT 704.900 1.400 705.740 614.600 ;
    RECT 706.020 1.400 706.860 614.600 ;
    RECT 707.140 1.400 707.980 614.600 ;
    RECT 708.260 1.400 709.100 614.600 ;
    RECT 709.380 1.400 710.220 614.600 ;
    RECT 710.500 1.400 711.340 614.600 ;
    RECT 711.620 1.400 712.460 614.600 ;
    RECT 712.740 1.400 713.580 614.600 ;
    RECT 713.860 1.400 714.700 614.600 ;
    RECT 714.980 1.400 715.820 614.600 ;
    RECT 716.100 1.400 716.940 614.600 ;
    RECT 717.220 1.400 718.060 614.600 ;
    RECT 718.340 1.400 719.180 614.600 ;
    RECT 719.460 1.400 720.300 614.600 ;
    RECT 720.580 1.400 721.420 614.600 ;
    RECT 721.700 1.400 722.540 614.600 ;
    RECT 722.820 1.400 723.660 614.600 ;
    RECT 723.940 1.400 724.780 614.600 ;
    RECT 725.060 1.400 725.900 614.600 ;
    RECT 726.180 1.400 727.020 614.600 ;
    RECT 727.300 1.400 728.140 614.600 ;
    RECT 728.420 1.400 729.260 614.600 ;
    RECT 729.540 1.400 730.380 614.600 ;
    RECT 730.660 1.400 731.500 614.600 ;
    RECT 731.780 1.400 732.620 614.600 ;
    RECT 732.900 1.400 733.740 614.600 ;
    RECT 734.020 1.400 734.860 614.600 ;
    RECT 735.140 1.400 735.980 614.600 ;
    RECT 736.260 1.400 737.100 614.600 ;
    RECT 737.380 1.400 738.220 614.600 ;
    RECT 738.500 1.400 739.340 614.600 ;
    RECT 739.620 1.400 740.460 614.600 ;
    RECT 740.740 1.400 741.580 614.600 ;
    RECT 741.860 1.400 742.700 614.600 ;
    RECT 742.980 1.400 743.820 614.600 ;
    RECT 744.100 1.400 744.940 614.600 ;
    RECT 745.220 1.400 746.060 614.600 ;
    RECT 746.340 1.400 747.180 614.600 ;
    RECT 747.460 1.400 748.300 614.600 ;
    RECT 748.580 1.400 749.420 614.600 ;
    RECT 749.700 1.400 750.540 614.600 ;
    RECT 750.820 1.400 751.660 614.600 ;
    RECT 751.940 1.400 752.780 614.600 ;
    RECT 753.060 1.400 753.900 614.600 ;
    RECT 754.180 1.400 755.020 614.600 ;
    RECT 755.300 1.400 756.140 614.600 ;
    RECT 756.420 1.400 757.260 614.600 ;
    RECT 757.540 1.400 758.380 614.600 ;
    RECT 758.660 1.400 759.500 614.600 ;
    RECT 759.780 1.400 760.620 614.600 ;
    RECT 760.900 1.400 761.740 614.600 ;
    RECT 762.020 1.400 762.860 614.600 ;
    RECT 763.140 1.400 763.980 614.600 ;
    RECT 764.260 1.400 765.100 614.600 ;
    RECT 765.380 1.400 766.220 614.600 ;
    RECT 766.500 1.400 767.340 614.600 ;
    RECT 767.620 1.400 768.460 614.600 ;
    RECT 768.740 1.400 769.580 614.600 ;
    RECT 769.860 1.400 770.700 614.600 ;
    RECT 770.980 1.400 771.820 614.600 ;
    RECT 772.100 1.400 772.940 614.600 ;
    RECT 773.220 1.400 774.060 614.600 ;
    RECT 774.340 1.400 775.180 614.600 ;
    RECT 775.460 1.400 776.300 614.600 ;
    RECT 776.580 1.400 777.420 614.600 ;
    RECT 777.700 1.400 778.540 614.600 ;
    RECT 778.820 1.400 779.660 614.600 ;
    RECT 779.940 1.400 780.780 614.600 ;
    RECT 781.060 1.400 781.900 614.600 ;
    RECT 782.180 1.400 783.020 614.600 ;
    RECT 783.300 1.400 784.140 614.600 ;
    RECT 784.420 1.400 785.260 614.600 ;
    RECT 785.540 1.400 786.380 614.600 ;
    RECT 786.660 1.400 787.500 614.600 ;
    RECT 787.780 1.400 788.620 614.600 ;
    RECT 788.900 1.400 789.740 614.600 ;
    RECT 790.020 1.400 790.860 614.600 ;
    RECT 791.140 1.400 791.980 614.600 ;
    RECT 792.260 1.400 793.100 614.600 ;
    RECT 793.380 1.400 794.220 614.600 ;
    RECT 794.500 1.400 795.340 614.600 ;
    RECT 795.620 1.400 796.460 614.600 ;
    RECT 796.740 1.400 797.580 614.600 ;
    RECT 797.860 1.400 798.700 614.600 ;
    RECT 798.980 1.400 799.820 614.600 ;
    RECT 800.100 1.400 800.940 614.600 ;
    RECT 801.220 1.400 802.060 614.600 ;
    RECT 802.340 1.400 803.180 614.600 ;
    RECT 803.460 1.400 804.300 614.600 ;
    RECT 804.580 1.400 805.420 614.600 ;
    RECT 805.700 1.400 806.540 614.600 ;
    RECT 806.820 1.400 807.660 614.600 ;
    RECT 807.940 1.400 808.780 614.600 ;
    RECT 809.060 1.400 809.900 614.600 ;
    RECT 810.180 1.400 811.020 614.600 ;
    RECT 811.300 1.400 812.140 614.600 ;
    RECT 812.420 1.400 813.260 614.600 ;
    RECT 813.540 1.400 814.380 614.600 ;
    RECT 814.660 1.400 815.500 614.600 ;
    RECT 815.780 1.400 816.620 614.600 ;
    RECT 816.900 1.400 817.740 614.600 ;
    RECT 818.020 1.400 818.860 614.600 ;
    RECT 819.140 1.400 819.980 614.600 ;
    RECT 820.260 1.400 821.100 614.600 ;
    RECT 821.380 1.400 822.220 614.600 ;
    RECT 822.500 1.400 823.340 614.600 ;
    RECT 823.620 1.400 824.460 614.600 ;
    RECT 824.740 1.400 825.580 614.600 ;
    RECT 825.860 1.400 826.700 614.600 ;
    RECT 826.980 1.400 827.820 614.600 ;
    RECT 828.100 1.400 828.940 614.600 ;
    RECT 829.220 1.400 830.060 614.600 ;
    RECT 830.340 1.400 831.180 614.600 ;
    RECT 831.460 1.400 832.300 614.600 ;
    RECT 832.580 1.400 833.420 614.600 ;
    RECT 833.700 1.400 834.540 614.600 ;
    RECT 834.820 1.400 835.660 614.600 ;
    RECT 835.940 1.400 836.780 614.600 ;
    RECT 837.060 1.400 837.900 614.600 ;
    RECT 838.180 1.400 839.020 614.600 ;
    RECT 839.300 1.400 840.140 614.600 ;
    RECT 840.420 1.400 841.260 614.600 ;
    RECT 841.540 1.400 842.380 614.600 ;
    RECT 842.660 1.400 843.500 614.600 ;
    RECT 843.780 1.400 844.620 614.600 ;
    RECT 844.900 1.400 845.740 614.600 ;
    RECT 846.020 1.400 846.860 614.600 ;
    RECT 847.140 1.400 847.980 614.600 ;
    RECT 848.260 1.400 849.100 614.600 ;
    RECT 849.380 1.400 850.220 614.600 ;
    RECT 850.500 1.400 851.340 614.600 ;
    RECT 851.620 1.400 852.460 614.600 ;
    RECT 852.740 1.400 853.580 614.600 ;
    RECT 853.860 1.400 854.700 614.600 ;
    RECT 854.980 1.400 855.820 614.600 ;
    RECT 856.100 1.400 856.940 614.600 ;
    RECT 857.220 1.400 858.060 614.600 ;
    RECT 858.340 1.400 859.180 614.600 ;
    RECT 859.460 1.400 860.300 614.600 ;
    RECT 860.580 1.400 861.420 614.600 ;
    RECT 861.700 1.400 862.540 614.600 ;
    RECT 862.820 1.400 863.660 614.600 ;
    RECT 863.940 1.400 864.780 614.600 ;
    RECT 865.060 1.400 865.900 614.600 ;
    RECT 866.180 1.400 867.020 614.600 ;
    RECT 867.300 1.400 868.140 614.600 ;
    RECT 868.420 1.400 869.260 614.600 ;
    RECT 869.540 1.400 870.380 614.600 ;
    RECT 870.660 1.400 871.500 614.600 ;
    RECT 871.780 1.400 872.620 614.600 ;
    RECT 872.900 1.400 873.740 614.600 ;
    RECT 874.020 1.400 874.860 614.600 ;
    RECT 875.140 1.400 875.980 614.600 ;
    RECT 876.260 1.400 877.100 614.600 ;
    RECT 877.380 1.400 878.220 614.600 ;
    RECT 878.500 1.400 879.340 614.600 ;
    RECT 879.620 1.400 880.460 614.600 ;
    RECT 880.740 1.400 881.580 614.600 ;
    RECT 881.860 1.400 882.700 614.600 ;
    RECT 882.980 1.400 883.820 614.600 ;
    RECT 884.100 1.400 884.940 614.600 ;
    RECT 885.220 1.400 886.060 614.600 ;
    RECT 886.340 1.400 887.180 614.600 ;
    RECT 887.460 1.400 888.300 614.600 ;
    RECT 888.580 1.400 889.420 614.600 ;
    RECT 889.700 1.400 890.540 614.600 ;
    RECT 890.820 1.400 891.660 614.600 ;
    RECT 891.940 1.400 892.780 614.600 ;
    RECT 893.060 1.400 893.900 614.600 ;
    RECT 894.180 1.400 895.020 614.600 ;
    RECT 895.300 1.400 896.140 614.600 ;
    RECT 896.420 1.400 897.260 614.600 ;
    RECT 897.540 1.400 898.380 614.600 ;
    RECT 898.660 1.400 899.500 614.600 ;
    RECT 899.780 1.400 900.620 614.600 ;
    RECT 900.900 1.400 901.740 614.600 ;
    RECT 902.020 1.400 902.860 614.600 ;
    RECT 903.140 1.400 903.980 614.600 ;
    RECT 904.260 1.400 905.100 614.600 ;
    RECT 905.380 1.400 906.220 614.600 ;
    RECT 906.500 1.400 907.340 614.600 ;
    RECT 907.620 1.400 908.460 614.600 ;
    RECT 908.740 1.400 909.580 614.600 ;
    RECT 909.860 1.400 910.700 614.600 ;
    RECT 910.980 1.400 911.820 614.600 ;
    RECT 912.100 1.400 912.940 614.600 ;
    RECT 913.220 1.400 914.060 614.600 ;
    RECT 914.340 1.400 915.180 614.600 ;
    RECT 915.460 1.400 916.300 614.600 ;
    RECT 916.580 1.400 917.420 614.600 ;
    RECT 917.700 1.400 918.540 614.600 ;
    RECT 918.820 1.400 919.660 614.600 ;
    RECT 919.940 1.400 920.780 614.600 ;
    RECT 921.060 1.400 921.900 614.600 ;
    RECT 922.180 1.400 923.020 614.600 ;
    RECT 923.300 1.400 924.140 614.600 ;
    RECT 924.420 1.400 925.260 614.600 ;
    RECT 925.540 1.400 926.380 614.600 ;
    RECT 926.660 1.400 927.500 614.600 ;
    RECT 927.780 1.400 928.620 614.600 ;
    RECT 928.900 1.400 929.740 614.600 ;
    RECT 930.020 1.400 930.860 614.600 ;
    RECT 931.140 1.400 931.980 614.600 ;
    RECT 932.260 1.400 933.100 614.600 ;
    RECT 933.380 1.400 934.220 614.600 ;
    RECT 934.500 1.400 935.340 614.600 ;
    RECT 935.620 1.400 936.460 614.600 ;
    RECT 936.740 1.400 937.580 614.600 ;
    RECT 937.860 1.400 938.700 614.600 ;
    RECT 938.980 1.400 939.820 614.600 ;
    RECT 940.100 1.400 940.940 614.600 ;
    RECT 941.220 1.400 942.060 614.600 ;
    RECT 942.340 1.400 943.180 614.600 ;
    RECT 943.460 1.400 944.300 614.600 ;
    RECT 944.580 1.400 945.420 614.600 ;
    RECT 945.700 1.400 946.540 614.600 ;
    RECT 946.820 1.400 947.660 614.600 ;
    RECT 947.940 1.400 948.780 614.600 ;
    RECT 949.060 1.400 949.900 614.600 ;
    RECT 950.180 1.400 951.020 614.600 ;
    RECT 951.300 1.400 952.140 614.600 ;
    RECT 952.420 1.400 953.260 614.600 ;
    RECT 953.540 1.400 954.380 614.600 ;
    RECT 954.660 1.400 955.500 614.600 ;
    RECT 955.780 1.400 956.620 614.600 ;
    RECT 956.900 1.400 957.740 614.600 ;
    RECT 958.020 1.400 958.860 614.600 ;
    RECT 959.140 1.400 959.980 614.600 ;
    RECT 960.260 1.400 961.100 614.600 ;
    RECT 961.380 1.400 962.220 614.600 ;
    RECT 962.500 1.400 963.340 614.600 ;
    RECT 963.620 1.400 964.460 614.600 ;
    RECT 964.740 1.400 965.580 614.600 ;
    RECT 965.860 1.400 966.700 614.600 ;
    RECT 966.980 1.400 967.820 614.600 ;
    RECT 968.100 1.400 968.940 614.600 ;
    RECT 969.220 1.400 970.060 614.600 ;
    RECT 970.340 1.400 971.180 614.600 ;
    RECT 971.460 1.400 972.300 614.600 ;
    RECT 972.580 1.400 973.420 614.600 ;
    RECT 973.700 1.400 974.540 614.600 ;
    RECT 974.820 1.400 975.660 614.600 ;
    RECT 975.940 1.400 976.780 614.600 ;
    RECT 977.060 1.400 977.900 614.600 ;
    RECT 978.180 1.400 979.020 614.600 ;
    RECT 979.300 1.400 980.140 614.600 ;
    RECT 980.420 1.400 981.260 614.600 ;
    RECT 981.540 1.400 982.380 614.600 ;
    RECT 982.660 1.400 983.500 614.600 ;
    RECT 983.780 1.400 984.620 614.600 ;
    RECT 984.900 1.400 985.740 614.600 ;
    RECT 986.020 1.400 986.860 614.600 ;
    RECT 987.140 1.400 987.980 614.600 ;
    RECT 988.260 1.400 989.100 614.600 ;
    RECT 989.380 1.400 990.220 614.600 ;
    RECT 990.500 1.400 991.340 614.600 ;
    RECT 991.620 1.400 992.460 614.600 ;
    RECT 992.740 1.400 993.580 614.600 ;
    RECT 993.860 1.400 994.700 614.600 ;
    RECT 994.980 1.400 995.820 614.600 ;
    RECT 996.100 1.400 996.940 614.600 ;
    RECT 997.220 1.400 998.060 614.600 ;
    RECT 998.340 1.400 999.180 614.600 ;
    RECT 999.460 1.400 1000.300 614.600 ;
    RECT 1000.580 1.400 1001.420 614.600 ;
    RECT 1001.700 1.400 1002.540 614.600 ;
    RECT 1002.820 1.400 1003.660 614.600 ;
    RECT 1003.940 1.400 1004.780 614.600 ;
    RECT 1005.060 1.400 1005.900 614.600 ;
    RECT 1006.180 1.400 1007.020 614.600 ;
    RECT 1007.300 1.400 1008.140 614.600 ;
    RECT 1008.420 1.400 1010.230 614.600 ;
    LAYER OVERLAP ;
    RECT 0 0 1010.230 616.000 ;
  END
END sram_32x16384_1rw

END LIBRARY
