VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_2848x32_1rw
  FOREIGN sram_2848x32_1rw 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 2078.600 BY 1618.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.505 0.070 1.575 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.645 0.070 1.715 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.785 0.070 1.855 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.925 0.070 1.995 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.345 0.070 2.415 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.625 0.070 2.695 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.185 0.070 3.255 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.025 0.070 4.095 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.445 0.070 4.515 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.865 0.070 4.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.145 0.070 5.215 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.705 0.070 5.775 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.125 0.070 6.195 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.545 0.070 6.615 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.825 0.070 6.895 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.385 0.070 7.455 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.225 0.070 8.295 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.505 0.070 8.575 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.065 0.070 9.135 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.345 0.070 9.415 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.485 0.070 9.555 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.905 0.070 9.975 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.745 0.070 10.815 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.025 0.070 11.095 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.585 0.070 11.655 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.425 0.070 12.495 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.705 0.070 12.775 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.265 0.070 13.335 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.545 0.070 13.615 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.105 0.070 14.175 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.385 0.070 14.455 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.525 0.070 14.595 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.945 0.070 15.015 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.225 0.070 15.295 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.645 0.070 15.715 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.785 0.070 15.855 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.205 0.070 16.275 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.625 0.070 16.695 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.905 0.070 16.975 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.465 0.070 17.535 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.745 0.070 17.815 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.885 0.070 17.955 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.305 0.070 18.375 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.585 0.070 18.655 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.725 0.070 18.795 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.145 0.070 19.215 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.425 0.070 19.495 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.985 0.070 20.055 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.685 0.070 20.755 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.825 0.070 20.895 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.105 0.070 21.175 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.245 0.070 21.315 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[143]
  PIN w_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[144]
  PIN w_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.665 0.070 21.735 ;
    END
  END w_mask_in[145]
  PIN w_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[146]
  PIN w_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END w_mask_in[147]
  PIN w_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.085 0.070 22.155 ;
    END
  END w_mask_in[148]
  PIN w_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[149]
  PIN w_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[150]
  PIN w_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.505 0.070 22.575 ;
    END
  END w_mask_in[151]
  PIN w_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[152]
  PIN w_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.785 0.070 22.855 ;
    END
  END w_mask_in[153]
  PIN w_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[154]
  PIN w_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[155]
  PIN w_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[156]
  PIN w_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.345 0.070 23.415 ;
    END
  END w_mask_in[157]
  PIN w_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[158]
  PIN w_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.625 0.070 23.695 ;
    END
  END w_mask_in[159]
  PIN w_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[160]
  PIN w_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[161]
  PIN w_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END w_mask_in[162]
  PIN w_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.185 0.070 24.255 ;
    END
  END w_mask_in[163]
  PIN w_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[164]
  PIN w_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END w_mask_in[165]
  PIN w_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.605 0.070 24.675 ;
    END
  END w_mask_in[166]
  PIN w_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[167]
  PIN w_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[168]
  PIN w_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.025 0.070 25.095 ;
    END
  END w_mask_in[169]
  PIN w_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[170]
  PIN w_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.305 0.070 25.375 ;
    END
  END w_mask_in[171]
  PIN w_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END w_mask_in[172]
  PIN w_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[173]
  PIN w_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.725 0.070 25.795 ;
    END
  END w_mask_in[174]
  PIN w_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END w_mask_in[175]
  PIN w_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[176]
  PIN w_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.145 0.070 26.215 ;
    END
  END w_mask_in[177]
  PIN w_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.285 0.070 26.355 ;
    END
  END w_mask_in[178]
  PIN w_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END w_mask_in[179]
  PIN w_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[180]
  PIN w_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.705 0.070 26.775 ;
    END
  END w_mask_in[181]
  PIN w_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[182]
  PIN w_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.985 0.070 27.055 ;
    END
  END w_mask_in[183]
  PIN w_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.125 0.070 27.195 ;
    END
  END w_mask_in[184]
  PIN w_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[185]
  PIN w_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.405 0.070 27.475 ;
    END
  END w_mask_in[186]
  PIN w_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.545 0.070 27.615 ;
    END
  END w_mask_in[187]
  PIN w_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[188]
  PIN w_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_in[189]
  PIN w_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[190]
  PIN w_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END w_mask_in[191]
  PIN w_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END w_mask_in[192]
  PIN w_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.385 0.070 28.455 ;
    END
  END w_mask_in[193]
  PIN w_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[194]
  PIN w_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.665 0.070 28.735 ;
    END
  END w_mask_in[195]
  PIN w_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END w_mask_in[196]
  PIN w_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.945 0.070 29.015 ;
    END
  END w_mask_in[197]
  PIN w_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END w_mask_in[198]
  PIN w_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.225 0.070 29.295 ;
    END
  END w_mask_in[199]
  PIN w_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[200]
  PIN w_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.505 0.070 29.575 ;
    END
  END w_mask_in[201]
  PIN w_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.645 0.070 29.715 ;
    END
  END w_mask_in[202]
  PIN w_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END w_mask_in[203]
  PIN w_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END w_mask_in[204]
  PIN w_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.065 0.070 30.135 ;
    END
  END w_mask_in[205]
  PIN w_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END w_mask_in[206]
  PIN w_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.345 0.070 30.415 ;
    END
  END w_mask_in[207]
  PIN w_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END w_mask_in[208]
  PIN w_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END w_mask_in[209]
  PIN w_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[210]
  PIN w_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.905 0.070 30.975 ;
    END
  END w_mask_in[211]
  PIN w_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END w_mask_in[212]
  PIN w_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.185 0.070 31.255 ;
    END
  END w_mask_in[213]
  PIN w_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.325 0.070 31.395 ;
    END
  END w_mask_in[214]
  PIN w_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[215]
  PIN w_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END w_mask_in[216]
  PIN w_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.745 0.070 31.815 ;
    END
  END w_mask_in[217]
  PIN w_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END w_mask_in[218]
  PIN w_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.025 0.070 32.095 ;
    END
  END w_mask_in[219]
  PIN w_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[220]
  PIN w_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END w_mask_in[221]
  PIN w_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END w_mask_in[222]
  PIN w_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.585 0.070 32.655 ;
    END
  END w_mask_in[223]
  PIN w_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END w_mask_in[224]
  PIN w_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.865 0.070 32.935 ;
    END
  END w_mask_in[225]
  PIN w_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.005 0.070 33.075 ;
    END
  END w_mask_in[226]
  PIN w_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END w_mask_in[227]
  PIN w_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[228]
  PIN w_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.425 0.070 33.495 ;
    END
  END w_mask_in[229]
  PIN w_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[230]
  PIN w_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_in[231]
  PIN w_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.845 0.070 33.915 ;
    END
  END w_mask_in[232]
  PIN w_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.985 0.070 34.055 ;
    END
  END w_mask_in[233]
  PIN w_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_in[234]
  PIN w_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.265 0.070 34.335 ;
    END
  END w_mask_in[235]
  PIN w_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[236]
  PIN w_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.545 0.070 34.615 ;
    END
  END w_mask_in[237]
  PIN w_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.685 0.070 34.755 ;
    END
  END w_mask_in[238]
  PIN w_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END w_mask_in[239]
  PIN w_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[240]
  PIN w_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.105 0.070 35.175 ;
    END
  END w_mask_in[241]
  PIN w_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END w_mask_in[242]
  PIN w_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.385 0.070 35.455 ;
    END
  END w_mask_in[243]
  PIN w_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.525 0.070 35.595 ;
    END
  END w_mask_in[244]
  PIN w_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END w_mask_in[245]
  PIN w_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END w_mask_in[246]
  PIN w_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.945 0.070 36.015 ;
    END
  END w_mask_in[247]
  PIN w_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END w_mask_in[248]
  PIN w_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.225 0.070 36.295 ;
    END
  END w_mask_in[249]
  PIN w_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.365 0.070 36.435 ;
    END
  END w_mask_in[250]
  PIN w_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END w_mask_in[251]
  PIN w_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[252]
  PIN w_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.785 0.070 36.855 ;
    END
  END w_mask_in[253]
  PIN w_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END w_mask_in[254]
  PIN w_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END w_mask_in[255]
  PIN w_mask_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.205 0.070 37.275 ;
    END
  END w_mask_in[256]
  PIN w_mask_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END w_mask_in[257]
  PIN w_mask_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END w_mask_in[258]
  PIN w_mask_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.625 0.070 37.695 ;
    END
  END w_mask_in[259]
  PIN w_mask_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[260]
  PIN w_mask_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.905 0.070 37.975 ;
    END
  END w_mask_in[261]
  PIN w_mask_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.045 0.070 38.115 ;
    END
  END w_mask_in[262]
  PIN w_mask_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END w_mask_in[263]
  PIN w_mask_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END w_mask_in[264]
  PIN w_mask_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.465 0.070 38.535 ;
    END
  END w_mask_in[265]
  PIN w_mask_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_in[266]
  PIN w_mask_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.745 0.070 38.815 ;
    END
  END w_mask_in[267]
  PIN w_mask_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.885 0.070 38.955 ;
    END
  END w_mask_in[268]
  PIN w_mask_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END w_mask_in[269]
  PIN w_mask_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[270]
  PIN w_mask_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.305 0.070 39.375 ;
    END
  END w_mask_in[271]
  PIN w_mask_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END w_mask_in[272]
  PIN w_mask_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END w_mask_in[273]
  PIN w_mask_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.725 0.070 39.795 ;
    END
  END w_mask_in[274]
  PIN w_mask_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END w_mask_in[275]
  PIN w_mask_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END w_mask_in[276]
  PIN w_mask_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.145 0.070 40.215 ;
    END
  END w_mask_in[277]
  PIN w_mask_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_in[278]
  PIN w_mask_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.425 0.070 40.495 ;
    END
  END w_mask_in[279]
  PIN w_mask_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[280]
  PIN w_mask_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END w_mask_in[281]
  PIN w_mask_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END w_mask_in[282]
  PIN w_mask_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.985 0.070 41.055 ;
    END
  END w_mask_in[283]
  PIN w_mask_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END w_mask_in[284]
  PIN w_mask_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END w_mask_in[285]
  PIN w_mask_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.405 0.070 41.475 ;
    END
  END w_mask_in[286]
  PIN w_mask_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END w_mask_in[287]
  PIN w_mask_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END w_mask_in[288]
  PIN w_mask_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.825 0.070 41.895 ;
    END
  END w_mask_in[289]
  PIN w_mask_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_in[290]
  PIN w_mask_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.105 0.070 42.175 ;
    END
  END w_mask_in[291]
  PIN w_mask_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.245 0.070 42.315 ;
    END
  END w_mask_in[292]
  PIN w_mask_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END w_mask_in[293]
  PIN w_mask_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_in[294]
  PIN w_mask_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.665 0.070 42.735 ;
    END
  END w_mask_in[295]
  PIN w_mask_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END w_mask_in[296]
  PIN w_mask_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END w_mask_in[297]
  PIN w_mask_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.085 0.070 43.155 ;
    END
  END w_mask_in[298]
  PIN w_mask_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END w_mask_in[299]
  PIN w_mask_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[300]
  PIN w_mask_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.505 0.070 43.575 ;
    END
  END w_mask_in[301]
  PIN w_mask_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END w_mask_in[302]
  PIN w_mask_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.785 0.070 43.855 ;
    END
  END w_mask_in[303]
  PIN w_mask_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END w_mask_in[304]
  PIN w_mask_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END w_mask_in[305]
  PIN w_mask_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END w_mask_in[306]
  PIN w_mask_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.345 0.070 44.415 ;
    END
  END w_mask_in[307]
  PIN w_mask_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END w_mask_in[308]
  PIN w_mask_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.625 0.070 44.695 ;
    END
  END w_mask_in[309]
  PIN w_mask_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END w_mask_in[310]
  PIN w_mask_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END w_mask_in[311]
  PIN w_mask_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END w_mask_in[312]
  PIN w_mask_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.185 0.070 45.255 ;
    END
  END w_mask_in[313]
  PIN w_mask_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END w_mask_in[314]
  PIN w_mask_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_in[315]
  PIN w_mask_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.605 0.070 45.675 ;
    END
  END w_mask_in[316]
  PIN w_mask_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END w_mask_in[317]
  PIN w_mask_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END w_mask_in[318]
  PIN w_mask_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.025 0.070 46.095 ;
    END
  END w_mask_in[319]
  PIN w_mask_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[320]
  PIN w_mask_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.305 0.070 46.375 ;
    END
  END w_mask_in[321]
  PIN w_mask_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END w_mask_in[322]
  PIN w_mask_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END w_mask_in[323]
  PIN w_mask_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END w_mask_in[324]
  PIN w_mask_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END w_mask_in[325]
  PIN w_mask_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END w_mask_in[326]
  PIN w_mask_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END w_mask_in[327]
  PIN w_mask_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.285 0.070 47.355 ;
    END
  END w_mask_in[328]
  PIN w_mask_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END w_mask_in[329]
  PIN w_mask_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_in[330]
  PIN w_mask_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.705 0.070 47.775 ;
    END
  END w_mask_in[331]
  PIN w_mask_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END w_mask_in[332]
  PIN w_mask_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.985 0.070 48.055 ;
    END
  END w_mask_in[333]
  PIN w_mask_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.125 0.070 48.195 ;
    END
  END w_mask_in[334]
  PIN w_mask_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END w_mask_in[335]
  PIN w_mask_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_in[336]
  PIN w_mask_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.545 0.070 48.615 ;
    END
  END w_mask_in[337]
  PIN w_mask_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END w_mask_in[338]
  PIN w_mask_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.825 0.070 48.895 ;
    END
  END w_mask_in[339]
  PIN w_mask_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END w_mask_in[340]
  PIN w_mask_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END w_mask_in[341]
  PIN w_mask_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END w_mask_in[342]
  PIN w_mask_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.385 0.070 49.455 ;
    END
  END w_mask_in[343]
  PIN w_mask_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END w_mask_in[344]
  PIN w_mask_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.665 0.070 49.735 ;
    END
  END w_mask_in[345]
  PIN w_mask_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.805 0.070 49.875 ;
    END
  END w_mask_in[346]
  PIN w_mask_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END w_mask_in[347]
  PIN w_mask_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.085 0.070 50.155 ;
    END
  END w_mask_in[348]
  PIN w_mask_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.225 0.070 50.295 ;
    END
  END w_mask_in[349]
  PIN w_mask_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_in[350]
  PIN w_mask_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.505 0.070 50.575 ;
    END
  END w_mask_in[351]
  PIN w_mask_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.645 0.070 50.715 ;
    END
  END w_mask_in[352]
  PIN w_mask_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END w_mask_in[353]
  PIN w_mask_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.925 0.070 50.995 ;
    END
  END w_mask_in[354]
  PIN w_mask_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.065 0.070 51.135 ;
    END
  END w_mask_in[355]
  PIN w_mask_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END w_mask_in[356]
  PIN w_mask_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.345 0.070 51.415 ;
    END
  END w_mask_in[357]
  PIN w_mask_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.485 0.070 51.555 ;
    END
  END w_mask_in[358]
  PIN w_mask_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END w_mask_in[359]
  PIN w_mask_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[360]
  PIN w_mask_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.905 0.070 51.975 ;
    END
  END w_mask_in[361]
  PIN w_mask_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END w_mask_in[362]
  PIN w_mask_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.185 0.070 52.255 ;
    END
  END w_mask_in[363]
  PIN w_mask_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END w_mask_in[364]
  PIN w_mask_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END w_mask_in[365]
  PIN w_mask_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.605 0.070 52.675 ;
    END
  END w_mask_in[366]
  PIN w_mask_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.745 0.070 52.815 ;
    END
  END w_mask_in[367]
  PIN w_mask_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END w_mask_in[368]
  PIN w_mask_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.025 0.070 53.095 ;
    END
  END w_mask_in[369]
  PIN w_mask_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.165 0.070 53.235 ;
    END
  END w_mask_in[370]
  PIN w_mask_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END w_mask_in[371]
  PIN w_mask_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.445 0.070 53.515 ;
    END
  END w_mask_in[372]
  PIN w_mask_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.585 0.070 53.655 ;
    END
  END w_mask_in[373]
  PIN w_mask_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END w_mask_in[374]
  PIN w_mask_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.865 0.070 53.935 ;
    END
  END w_mask_in[375]
  PIN w_mask_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.005 0.070 54.075 ;
    END
  END w_mask_in[376]
  PIN w_mask_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END w_mask_in[377]
  PIN w_mask_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_in[378]
  PIN w_mask_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.425 0.070 54.495 ;
    END
  END w_mask_in[379]
  PIN w_mask_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[380]
  PIN w_mask_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.705 0.070 54.775 ;
    END
  END w_mask_in[381]
  PIN w_mask_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.845 0.070 54.915 ;
    END
  END w_mask_in[382]
  PIN w_mask_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END w_mask_in[383]
  PIN w_mask_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END w_mask_in[384]
  PIN w_mask_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.265 0.070 55.335 ;
    END
  END w_mask_in[385]
  PIN w_mask_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END w_mask_in[386]
  PIN w_mask_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.545 0.070 55.615 ;
    END
  END w_mask_in[387]
  PIN w_mask_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.685 0.070 55.755 ;
    END
  END w_mask_in[388]
  PIN w_mask_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END w_mask_in[389]
  PIN w_mask_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_in[390]
  PIN w_mask_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.105 0.070 56.175 ;
    END
  END w_mask_in[391]
  PIN w_mask_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END w_mask_in[392]
  PIN w_mask_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.385 0.070 56.455 ;
    END
  END w_mask_in[393]
  PIN w_mask_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.525 0.070 56.595 ;
    END
  END w_mask_in[394]
  PIN w_mask_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END w_mask_in[395]
  PIN w_mask_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END w_mask_in[396]
  PIN w_mask_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.945 0.070 57.015 ;
    END
  END w_mask_in[397]
  PIN w_mask_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END w_mask_in[398]
  PIN w_mask_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.225 0.070 57.295 ;
    END
  END w_mask_in[399]
  PIN w_mask_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END w_mask_in[400]
  PIN w_mask_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END w_mask_in[401]
  PIN w_mask_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END w_mask_in[402]
  PIN w_mask_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.785 0.070 57.855 ;
    END
  END w_mask_in[403]
  PIN w_mask_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END w_mask_in[404]
  PIN w_mask_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.065 0.070 58.135 ;
    END
  END w_mask_in[405]
  PIN w_mask_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END w_mask_in[406]
  PIN w_mask_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END w_mask_in[407]
  PIN w_mask_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END w_mask_in[408]
  PIN w_mask_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.625 0.070 58.695 ;
    END
  END w_mask_in[409]
  PIN w_mask_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END w_mask_in[410]
  PIN w_mask_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.905 0.070 58.975 ;
    END
  END w_mask_in[411]
  PIN w_mask_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.045 0.070 59.115 ;
    END
  END w_mask_in[412]
  PIN w_mask_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END w_mask_in[413]
  PIN w_mask_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.325 0.070 59.395 ;
    END
  END w_mask_in[414]
  PIN w_mask_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.465 0.070 59.535 ;
    END
  END w_mask_in[415]
  PIN w_mask_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END w_mask_in[416]
  PIN w_mask_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.745 0.070 59.815 ;
    END
  END w_mask_in[417]
  PIN w_mask_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END w_mask_in[418]
  PIN w_mask_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END w_mask_in[419]
  PIN w_mask_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[420]
  PIN w_mask_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.305 0.070 60.375 ;
    END
  END w_mask_in[421]
  PIN w_mask_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END w_mask_in[422]
  PIN w_mask_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.585 0.070 60.655 ;
    END
  END w_mask_in[423]
  PIN w_mask_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.725 0.070 60.795 ;
    END
  END w_mask_in[424]
  PIN w_mask_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END w_mask_in[425]
  PIN w_mask_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.005 0.070 61.075 ;
    END
  END w_mask_in[426]
  PIN w_mask_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.145 0.070 61.215 ;
    END
  END w_mask_in[427]
  PIN w_mask_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END w_mask_in[428]
  PIN w_mask_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.425 0.070 61.495 ;
    END
  END w_mask_in[429]
  PIN w_mask_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.565 0.070 61.635 ;
    END
  END w_mask_in[430]
  PIN w_mask_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END w_mask_in[431]
  PIN w_mask_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.845 0.070 61.915 ;
    END
  END w_mask_in[432]
  PIN w_mask_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.985 0.070 62.055 ;
    END
  END w_mask_in[433]
  PIN w_mask_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END w_mask_in[434]
  PIN w_mask_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.265 0.070 62.335 ;
    END
  END w_mask_in[435]
  PIN w_mask_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END w_mask_in[436]
  PIN w_mask_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END w_mask_in[437]
  PIN w_mask_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.685 0.070 62.755 ;
    END
  END w_mask_in[438]
  PIN w_mask_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.825 0.070 62.895 ;
    END
  END w_mask_in[439]
  PIN w_mask_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END w_mask_in[440]
  PIN w_mask_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.105 0.070 63.175 ;
    END
  END w_mask_in[441]
  PIN w_mask_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.245 0.070 63.315 ;
    END
  END w_mask_in[442]
  PIN w_mask_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END w_mask_in[443]
  PIN w_mask_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END w_mask_in[444]
  PIN w_mask_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.665 0.070 63.735 ;
    END
  END w_mask_in[445]
  PIN w_mask_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END w_mask_in[446]
  PIN w_mask_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.945 0.070 64.015 ;
    END
  END w_mask_in[447]
  PIN w_mask_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.085 0.070 64.155 ;
    END
  END w_mask_in[448]
  PIN w_mask_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END w_mask_in[449]
  PIN w_mask_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END w_mask_in[450]
  PIN w_mask_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.505 0.070 64.575 ;
    END
  END w_mask_in[451]
  PIN w_mask_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END w_mask_in[452]
  PIN w_mask_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.785 0.070 64.855 ;
    END
  END w_mask_in[453]
  PIN w_mask_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.925 0.070 64.995 ;
    END
  END w_mask_in[454]
  PIN w_mask_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END w_mask_in[455]
  PIN w_mask_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END w_mask_in[456]
  PIN w_mask_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.345 0.070 65.415 ;
    END
  END w_mask_in[457]
  PIN w_mask_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END w_mask_in[458]
  PIN w_mask_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.625 0.070 65.695 ;
    END
  END w_mask_in[459]
  PIN w_mask_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END w_mask_in[460]
  PIN w_mask_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.905 0.070 65.975 ;
    END
  END w_mask_in[461]
  PIN w_mask_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END w_mask_in[462]
  PIN w_mask_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.185 0.070 66.255 ;
    END
  END w_mask_in[463]
  PIN w_mask_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END w_mask_in[464]
  PIN w_mask_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.465 0.070 66.535 ;
    END
  END w_mask_in[465]
  PIN w_mask_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.605 0.070 66.675 ;
    END
  END w_mask_in[466]
  PIN w_mask_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END w_mask_in[467]
  PIN w_mask_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END w_mask_in[468]
  PIN w_mask_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.025 0.070 67.095 ;
    END
  END w_mask_in[469]
  PIN w_mask_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END w_mask_in[470]
  PIN w_mask_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.305 0.070 67.375 ;
    END
  END w_mask_in[471]
  PIN w_mask_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.445 0.070 67.515 ;
    END
  END w_mask_in[472]
  PIN w_mask_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END w_mask_in[473]
  PIN w_mask_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.725 0.070 67.795 ;
    END
  END w_mask_in[474]
  PIN w_mask_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.865 0.070 67.935 ;
    END
  END w_mask_in[475]
  PIN w_mask_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END w_mask_in[476]
  PIN w_mask_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.145 0.070 68.215 ;
    END
  END w_mask_in[477]
  PIN w_mask_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.285 0.070 68.355 ;
    END
  END w_mask_in[478]
  PIN w_mask_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END w_mask_in[479]
  PIN w_mask_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_in[480]
  PIN w_mask_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.705 0.070 68.775 ;
    END
  END w_mask_in[481]
  PIN w_mask_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END w_mask_in[482]
  PIN w_mask_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.985 0.070 69.055 ;
    END
  END w_mask_in[483]
  PIN w_mask_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END w_mask_in[484]
  PIN w_mask_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END w_mask_in[485]
  PIN w_mask_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.405 0.070 69.475 ;
    END
  END w_mask_in[486]
  PIN w_mask_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.545 0.070 69.615 ;
    END
  END w_mask_in[487]
  PIN w_mask_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END w_mask_in[488]
  PIN w_mask_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.825 0.070 69.895 ;
    END
  END w_mask_in[489]
  PIN w_mask_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END w_mask_in[490]
  PIN w_mask_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END w_mask_in[491]
  PIN w_mask_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END w_mask_in[492]
  PIN w_mask_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.385 0.070 70.455 ;
    END
  END w_mask_in[493]
  PIN w_mask_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END w_mask_in[494]
  PIN w_mask_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.665 0.070 70.735 ;
    END
  END w_mask_in[495]
  PIN w_mask_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END w_mask_in[496]
  PIN w_mask_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END w_mask_in[497]
  PIN w_mask_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END w_mask_in[498]
  PIN w_mask_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.225 0.070 71.295 ;
    END
  END w_mask_in[499]
  PIN w_mask_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END w_mask_in[500]
  PIN w_mask_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.505 0.070 71.575 ;
    END
  END w_mask_in[501]
  PIN w_mask_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.645 0.070 71.715 ;
    END
  END w_mask_in[502]
  PIN w_mask_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END w_mask_in[503]
  PIN w_mask_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END w_mask_in[504]
  PIN w_mask_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.065 0.070 72.135 ;
    END
  END w_mask_in[505]
  PIN w_mask_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END w_mask_in[506]
  PIN w_mask_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.345 0.070 72.415 ;
    END
  END w_mask_in[507]
  PIN w_mask_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END w_mask_in[508]
  PIN w_mask_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END w_mask_in[509]
  PIN w_mask_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END w_mask_in[510]
  PIN w_mask_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.905 0.070 72.975 ;
    END
  END w_mask_in[511]
  PIN w_mask_in[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END w_mask_in[512]
  PIN w_mask_in[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.185 0.070 73.255 ;
    END
  END w_mask_in[513]
  PIN w_mask_in[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.325 0.070 73.395 ;
    END
  END w_mask_in[514]
  PIN w_mask_in[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END w_mask_in[515]
  PIN w_mask_in[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END w_mask_in[516]
  PIN w_mask_in[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.745 0.070 73.815 ;
    END
  END w_mask_in[517]
  PIN w_mask_in[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END w_mask_in[518]
  PIN w_mask_in[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.025 0.070 74.095 ;
    END
  END w_mask_in[519]
  PIN w_mask_in[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END w_mask_in[520]
  PIN w_mask_in[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END w_mask_in[521]
  PIN w_mask_in[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.445 0.070 74.515 ;
    END
  END w_mask_in[522]
  PIN w_mask_in[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.585 0.070 74.655 ;
    END
  END w_mask_in[523]
  PIN w_mask_in[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END w_mask_in[524]
  PIN w_mask_in[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.865 0.070 74.935 ;
    END
  END w_mask_in[525]
  PIN w_mask_in[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END w_mask_in[526]
  PIN w_mask_in[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END w_mask_in[527]
  PIN w_mask_in[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END w_mask_in[528]
  PIN w_mask_in[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.425 0.070 75.495 ;
    END
  END w_mask_in[529]
  PIN w_mask_in[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END w_mask_in[530]
  PIN w_mask_in[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.705 0.070 75.775 ;
    END
  END w_mask_in[531]
  PIN w_mask_in[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END w_mask_in[532]
  PIN w_mask_in[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END w_mask_in[533]
  PIN w_mask_in[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.125 0.070 76.195 ;
    END
  END w_mask_in[534]
  PIN w_mask_in[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.265 0.070 76.335 ;
    END
  END w_mask_in[535]
  PIN w_mask_in[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END w_mask_in[536]
  PIN w_mask_in[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.545 0.070 76.615 ;
    END
  END w_mask_in[537]
  PIN w_mask_in[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.685 0.070 76.755 ;
    END
  END w_mask_in[538]
  PIN w_mask_in[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END w_mask_in[539]
  PIN w_mask_in[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END w_mask_in[540]
  PIN w_mask_in[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.105 0.070 77.175 ;
    END
  END w_mask_in[541]
  PIN w_mask_in[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END w_mask_in[542]
  PIN w_mask_in[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.385 0.070 77.455 ;
    END
  END w_mask_in[543]
  PIN w_mask_in[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.525 0.070 77.595 ;
    END
  END w_mask_in[544]
  PIN w_mask_in[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END w_mask_in[545]
  PIN w_mask_in[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END w_mask_in[546]
  PIN w_mask_in[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.945 0.070 78.015 ;
    END
  END w_mask_in[547]
  PIN w_mask_in[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END w_mask_in[548]
  PIN w_mask_in[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.225 0.070 78.295 ;
    END
  END w_mask_in[549]
  PIN w_mask_in[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END w_mask_in[550]
  PIN w_mask_in[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END w_mask_in[551]
  PIN w_mask_in[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.645 0.070 78.715 ;
    END
  END w_mask_in[552]
  PIN w_mask_in[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.785 0.070 78.855 ;
    END
  END w_mask_in[553]
  PIN w_mask_in[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END w_mask_in[554]
  PIN w_mask_in[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.065 0.070 79.135 ;
    END
  END w_mask_in[555]
  PIN w_mask_in[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.205 0.070 79.275 ;
    END
  END w_mask_in[556]
  PIN w_mask_in[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END w_mask_in[557]
  PIN w_mask_in[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.485 0.070 79.555 ;
    END
  END w_mask_in[558]
  PIN w_mask_in[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.625 0.070 79.695 ;
    END
  END w_mask_in[559]
  PIN w_mask_in[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END w_mask_in[560]
  PIN w_mask_in[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.905 0.070 79.975 ;
    END
  END w_mask_in[561]
  PIN w_mask_in[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.045 0.070 80.115 ;
    END
  END w_mask_in[562]
  PIN w_mask_in[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END w_mask_in[563]
  PIN w_mask_in[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.325 0.070 80.395 ;
    END
  END w_mask_in[564]
  PIN w_mask_in[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.465 0.070 80.535 ;
    END
  END w_mask_in[565]
  PIN w_mask_in[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END w_mask_in[566]
  PIN w_mask_in[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.745 0.070 80.815 ;
    END
  END w_mask_in[567]
  PIN w_mask_in[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.885 0.070 80.955 ;
    END
  END w_mask_in[568]
  PIN w_mask_in[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END w_mask_in[569]
  PIN w_mask_in[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END w_mask_in[570]
  PIN w_mask_in[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.305 0.070 81.375 ;
    END
  END w_mask_in[571]
  PIN w_mask_in[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END w_mask_in[572]
  PIN w_mask_in[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.585 0.070 81.655 ;
    END
  END w_mask_in[573]
  PIN w_mask_in[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.725 0.070 81.795 ;
    END
  END w_mask_in[574]
  PIN w_mask_in[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END w_mask_in[575]
  PIN w_mask_in[576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.005 0.070 82.075 ;
    END
  END w_mask_in[576]
  PIN w_mask_in[577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.145 0.070 82.215 ;
    END
  END w_mask_in[577]
  PIN w_mask_in[578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END w_mask_in[578]
  PIN w_mask_in[579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.425 0.070 82.495 ;
    END
  END w_mask_in[579]
  PIN w_mask_in[580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END w_mask_in[580]
  PIN w_mask_in[581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END w_mask_in[581]
  PIN w_mask_in[582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.845 0.070 82.915 ;
    END
  END w_mask_in[582]
  PIN w_mask_in[583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.985 0.070 83.055 ;
    END
  END w_mask_in[583]
  PIN w_mask_in[584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END w_mask_in[584]
  PIN w_mask_in[585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.265 0.070 83.335 ;
    END
  END w_mask_in[585]
  PIN w_mask_in[586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.405 0.070 83.475 ;
    END
  END w_mask_in[586]
  PIN w_mask_in[587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END w_mask_in[587]
  PIN w_mask_in[588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END w_mask_in[588]
  PIN w_mask_in[589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.825 0.070 83.895 ;
    END
  END w_mask_in[589]
  PIN w_mask_in[590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END w_mask_in[590]
  PIN w_mask_in[591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.105 0.070 84.175 ;
    END
  END w_mask_in[591]
  PIN w_mask_in[592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.245 0.070 84.315 ;
    END
  END w_mask_in[592]
  PIN w_mask_in[593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END w_mask_in[593]
  PIN w_mask_in[594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END w_mask_in[594]
  PIN w_mask_in[595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.665 0.070 84.735 ;
    END
  END w_mask_in[595]
  PIN w_mask_in[596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END w_mask_in[596]
  PIN w_mask_in[597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.945 0.070 85.015 ;
    END
  END w_mask_in[597]
  PIN w_mask_in[598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.085 0.070 85.155 ;
    END
  END w_mask_in[598]
  PIN w_mask_in[599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END w_mask_in[599]
  PIN w_mask_in[600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END w_mask_in[600]
  PIN w_mask_in[601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.505 0.070 85.575 ;
    END
  END w_mask_in[601]
  PIN w_mask_in[602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END w_mask_in[602]
  PIN w_mask_in[603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.785 0.070 85.855 ;
    END
  END w_mask_in[603]
  PIN w_mask_in[604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.925 0.070 85.995 ;
    END
  END w_mask_in[604]
  PIN w_mask_in[605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END w_mask_in[605]
  PIN w_mask_in[606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.205 0.070 86.275 ;
    END
  END w_mask_in[606]
  PIN w_mask_in[607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.345 0.070 86.415 ;
    END
  END w_mask_in[607]
  PIN w_mask_in[608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END w_mask_in[608]
  PIN w_mask_in[609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.625 0.070 86.695 ;
    END
  END w_mask_in[609]
  PIN w_mask_in[610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END w_mask_in[610]
  PIN w_mask_in[611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END w_mask_in[611]
  PIN w_mask_in[612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.045 0.070 87.115 ;
    END
  END w_mask_in[612]
  PIN w_mask_in[613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.185 0.070 87.255 ;
    END
  END w_mask_in[613]
  PIN w_mask_in[614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END w_mask_in[614]
  PIN w_mask_in[615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.465 0.070 87.535 ;
    END
  END w_mask_in[615]
  PIN w_mask_in[616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.605 0.070 87.675 ;
    END
  END w_mask_in[616]
  PIN w_mask_in[617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END w_mask_in[617]
  PIN w_mask_in[618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.885 0.070 87.955 ;
    END
  END w_mask_in[618]
  PIN w_mask_in[619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.025 0.070 88.095 ;
    END
  END w_mask_in[619]
  PIN w_mask_in[620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END w_mask_in[620]
  PIN w_mask_in[621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.305 0.070 88.375 ;
    END
  END w_mask_in[621]
  PIN w_mask_in[622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.445 0.070 88.515 ;
    END
  END w_mask_in[622]
  PIN w_mask_in[623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END w_mask_in[623]
  PIN w_mask_in[624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.725 0.070 88.795 ;
    END
  END w_mask_in[624]
  PIN w_mask_in[625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.865 0.070 88.935 ;
    END
  END w_mask_in[625]
  PIN w_mask_in[626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END w_mask_in[626]
  PIN w_mask_in[627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.145 0.070 89.215 ;
    END
  END w_mask_in[627]
  PIN w_mask_in[628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.285 0.070 89.355 ;
    END
  END w_mask_in[628]
  PIN w_mask_in[629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.425 0.070 89.495 ;
    END
  END w_mask_in[629]
  PIN w_mask_in[630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END w_mask_in[630]
  PIN w_mask_in[631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.705 0.070 89.775 ;
    END
  END w_mask_in[631]
  PIN w_mask_in[632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END w_mask_in[632]
  PIN w_mask_in[633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.985 0.070 90.055 ;
    END
  END w_mask_in[633]
  PIN w_mask_in[634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.125 0.070 90.195 ;
    END
  END w_mask_in[634]
  PIN w_mask_in[635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END w_mask_in[635]
  PIN w_mask_in[636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.405 0.070 90.475 ;
    END
  END w_mask_in[636]
  PIN w_mask_in[637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.545 0.070 90.615 ;
    END
  END w_mask_in[637]
  PIN w_mask_in[638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END w_mask_in[638]
  PIN w_mask_in[639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.825 0.070 90.895 ;
    END
  END w_mask_in[639]
  PIN w_mask_in[640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.965 0.070 91.035 ;
    END
  END w_mask_in[640]
  PIN w_mask_in[641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.105 0.070 91.175 ;
    END
  END w_mask_in[641]
  PIN w_mask_in[642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.245 0.070 91.315 ;
    END
  END w_mask_in[642]
  PIN w_mask_in[643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.385 0.070 91.455 ;
    END
  END w_mask_in[643]
  PIN w_mask_in[644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END w_mask_in[644]
  PIN w_mask_in[645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.665 0.070 91.735 ;
    END
  END w_mask_in[645]
  PIN w_mask_in[646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.805 0.070 91.875 ;
    END
  END w_mask_in[646]
  PIN w_mask_in[647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.945 0.070 92.015 ;
    END
  END w_mask_in[647]
  PIN w_mask_in[648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.085 0.070 92.155 ;
    END
  END w_mask_in[648]
  PIN w_mask_in[649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.225 0.070 92.295 ;
    END
  END w_mask_in[649]
  PIN w_mask_in[650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END w_mask_in[650]
  PIN w_mask_in[651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.505 0.070 92.575 ;
    END
  END w_mask_in[651]
  PIN w_mask_in[652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.645 0.070 92.715 ;
    END
  END w_mask_in[652]
  PIN w_mask_in[653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.785 0.070 92.855 ;
    END
  END w_mask_in[653]
  PIN w_mask_in[654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.925 0.070 92.995 ;
    END
  END w_mask_in[654]
  PIN w_mask_in[655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.065 0.070 93.135 ;
    END
  END w_mask_in[655]
  PIN w_mask_in[656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END w_mask_in[656]
  PIN w_mask_in[657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.345 0.070 93.415 ;
    END
  END w_mask_in[657]
  PIN w_mask_in[658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.485 0.070 93.555 ;
    END
  END w_mask_in[658]
  PIN w_mask_in[659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.625 0.070 93.695 ;
    END
  END w_mask_in[659]
  PIN w_mask_in[660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.765 0.070 93.835 ;
    END
  END w_mask_in[660]
  PIN w_mask_in[661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.905 0.070 93.975 ;
    END
  END w_mask_in[661]
  PIN w_mask_in[662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END w_mask_in[662]
  PIN w_mask_in[663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.185 0.070 94.255 ;
    END
  END w_mask_in[663]
  PIN w_mask_in[664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.325 0.070 94.395 ;
    END
  END w_mask_in[664]
  PIN w_mask_in[665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END w_mask_in[665]
  PIN w_mask_in[666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.605 0.070 94.675 ;
    END
  END w_mask_in[666]
  PIN w_mask_in[667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.745 0.070 94.815 ;
    END
  END w_mask_in[667]
  PIN w_mask_in[668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END w_mask_in[668]
  PIN w_mask_in[669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.025 0.070 95.095 ;
    END
  END w_mask_in[669]
  PIN w_mask_in[670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.165 0.070 95.235 ;
    END
  END w_mask_in[670]
  PIN w_mask_in[671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.305 0.070 95.375 ;
    END
  END w_mask_in[671]
  PIN w_mask_in[672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END w_mask_in[672]
  PIN w_mask_in[673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.585 0.070 95.655 ;
    END
  END w_mask_in[673]
  PIN w_mask_in[674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.725 0.070 95.795 ;
    END
  END w_mask_in[674]
  PIN w_mask_in[675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.865 0.070 95.935 ;
    END
  END w_mask_in[675]
  PIN w_mask_in[676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.005 0.070 96.075 ;
    END
  END w_mask_in[676]
  PIN w_mask_in[677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.145 0.070 96.215 ;
    END
  END w_mask_in[677]
  PIN w_mask_in[678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.285 0.070 96.355 ;
    END
  END w_mask_in[678]
  PIN w_mask_in[679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.425 0.070 96.495 ;
    END
  END w_mask_in[679]
  PIN w_mask_in[680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END w_mask_in[680]
  PIN w_mask_in[681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.705 0.070 96.775 ;
    END
  END w_mask_in[681]
  PIN w_mask_in[682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.845 0.070 96.915 ;
    END
  END w_mask_in[682]
  PIN w_mask_in[683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.985 0.070 97.055 ;
    END
  END w_mask_in[683]
  PIN w_mask_in[684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.125 0.070 97.195 ;
    END
  END w_mask_in[684]
  PIN w_mask_in[685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.265 0.070 97.335 ;
    END
  END w_mask_in[685]
  PIN w_mask_in[686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END w_mask_in[686]
  PIN w_mask_in[687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.545 0.070 97.615 ;
    END
  END w_mask_in[687]
  PIN w_mask_in[688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.685 0.070 97.755 ;
    END
  END w_mask_in[688]
  PIN w_mask_in[689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.825 0.070 97.895 ;
    END
  END w_mask_in[689]
  PIN w_mask_in[690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.965 0.070 98.035 ;
    END
  END w_mask_in[690]
  PIN w_mask_in[691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.105 0.070 98.175 ;
    END
  END w_mask_in[691]
  PIN w_mask_in[692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.245 0.070 98.315 ;
    END
  END w_mask_in[692]
  PIN w_mask_in[693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.385 0.070 98.455 ;
    END
  END w_mask_in[693]
  PIN w_mask_in[694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.525 0.070 98.595 ;
    END
  END w_mask_in[694]
  PIN w_mask_in[695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.665 0.070 98.735 ;
    END
  END w_mask_in[695]
  PIN w_mask_in[696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.805 0.070 98.875 ;
    END
  END w_mask_in[696]
  PIN w_mask_in[697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.945 0.070 99.015 ;
    END
  END w_mask_in[697]
  PIN w_mask_in[698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.085 0.070 99.155 ;
    END
  END w_mask_in[698]
  PIN w_mask_in[699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.225 0.070 99.295 ;
    END
  END w_mask_in[699]
  PIN w_mask_in[700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.365 0.070 99.435 ;
    END
  END w_mask_in[700]
  PIN w_mask_in[701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.505 0.070 99.575 ;
    END
  END w_mask_in[701]
  PIN w_mask_in[702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END w_mask_in[702]
  PIN w_mask_in[703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.785 0.070 99.855 ;
    END
  END w_mask_in[703]
  PIN w_mask_in[704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.925 0.070 99.995 ;
    END
  END w_mask_in[704]
  PIN w_mask_in[705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.065 0.070 100.135 ;
    END
  END w_mask_in[705]
  PIN w_mask_in[706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.205 0.070 100.275 ;
    END
  END w_mask_in[706]
  PIN w_mask_in[707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END w_mask_in[707]
  PIN w_mask_in[708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.485 0.070 100.555 ;
    END
  END w_mask_in[708]
  PIN w_mask_in[709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.625 0.070 100.695 ;
    END
  END w_mask_in[709]
  PIN w_mask_in[710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END w_mask_in[710]
  PIN w_mask_in[711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.905 0.070 100.975 ;
    END
  END w_mask_in[711]
  PIN w_mask_in[712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.045 0.070 101.115 ;
    END
  END w_mask_in[712]
  PIN w_mask_in[713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.185 0.070 101.255 ;
    END
  END w_mask_in[713]
  PIN w_mask_in[714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END w_mask_in[714]
  PIN w_mask_in[715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.465 0.070 101.535 ;
    END
  END w_mask_in[715]
  PIN w_mask_in[716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END w_mask_in[716]
  PIN w_mask_in[717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.745 0.070 101.815 ;
    END
  END w_mask_in[717]
  PIN w_mask_in[718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.885 0.070 101.955 ;
    END
  END w_mask_in[718]
  PIN w_mask_in[719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.025 0.070 102.095 ;
    END
  END w_mask_in[719]
  PIN w_mask_in[720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.165 0.070 102.235 ;
    END
  END w_mask_in[720]
  PIN w_mask_in[721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.305 0.070 102.375 ;
    END
  END w_mask_in[721]
  PIN w_mask_in[722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END w_mask_in[722]
  PIN w_mask_in[723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.585 0.070 102.655 ;
    END
  END w_mask_in[723]
  PIN w_mask_in[724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.725 0.070 102.795 ;
    END
  END w_mask_in[724]
  PIN w_mask_in[725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.865 0.070 102.935 ;
    END
  END w_mask_in[725]
  PIN w_mask_in[726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.005 0.070 103.075 ;
    END
  END w_mask_in[726]
  PIN w_mask_in[727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.145 0.070 103.215 ;
    END
  END w_mask_in[727]
  PIN w_mask_in[728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END w_mask_in[728]
  PIN w_mask_in[729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.425 0.070 103.495 ;
    END
  END w_mask_in[729]
  PIN w_mask_in[730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.565 0.070 103.635 ;
    END
  END w_mask_in[730]
  PIN w_mask_in[731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.705 0.070 103.775 ;
    END
  END w_mask_in[731]
  PIN w_mask_in[732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.845 0.070 103.915 ;
    END
  END w_mask_in[732]
  PIN w_mask_in[733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.985 0.070 104.055 ;
    END
  END w_mask_in[733]
  PIN w_mask_in[734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.125 0.070 104.195 ;
    END
  END w_mask_in[734]
  PIN w_mask_in[735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.265 0.070 104.335 ;
    END
  END w_mask_in[735]
  PIN w_mask_in[736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.405 0.070 104.475 ;
    END
  END w_mask_in[736]
  PIN w_mask_in[737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.545 0.070 104.615 ;
    END
  END w_mask_in[737]
  PIN w_mask_in[738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.685 0.070 104.755 ;
    END
  END w_mask_in[738]
  PIN w_mask_in[739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.825 0.070 104.895 ;
    END
  END w_mask_in[739]
  PIN w_mask_in[740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.965 0.070 105.035 ;
    END
  END w_mask_in[740]
  PIN w_mask_in[741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.105 0.070 105.175 ;
    END
  END w_mask_in[741]
  PIN w_mask_in[742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END w_mask_in[742]
  PIN w_mask_in[743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.385 0.070 105.455 ;
    END
  END w_mask_in[743]
  PIN w_mask_in[744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.525 0.070 105.595 ;
    END
  END w_mask_in[744]
  PIN w_mask_in[745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.665 0.070 105.735 ;
    END
  END w_mask_in[745]
  PIN w_mask_in[746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END w_mask_in[746]
  PIN w_mask_in[747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.945 0.070 106.015 ;
    END
  END w_mask_in[747]
  PIN w_mask_in[748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.085 0.070 106.155 ;
    END
  END w_mask_in[748]
  PIN w_mask_in[749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.225 0.070 106.295 ;
    END
  END w_mask_in[749]
  PIN w_mask_in[750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.365 0.070 106.435 ;
    END
  END w_mask_in[750]
  PIN w_mask_in[751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.505 0.070 106.575 ;
    END
  END w_mask_in[751]
  PIN w_mask_in[752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.645 0.070 106.715 ;
    END
  END w_mask_in[752]
  PIN w_mask_in[753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.785 0.070 106.855 ;
    END
  END w_mask_in[753]
  PIN w_mask_in[754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.925 0.070 106.995 ;
    END
  END w_mask_in[754]
  PIN w_mask_in[755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.065 0.070 107.135 ;
    END
  END w_mask_in[755]
  PIN w_mask_in[756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END w_mask_in[756]
  PIN w_mask_in[757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.345 0.070 107.415 ;
    END
  END w_mask_in[757]
  PIN w_mask_in[758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END w_mask_in[758]
  PIN w_mask_in[759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.625 0.070 107.695 ;
    END
  END w_mask_in[759]
  PIN w_mask_in[760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.765 0.070 107.835 ;
    END
  END w_mask_in[760]
  PIN w_mask_in[761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.905 0.070 107.975 ;
    END
  END w_mask_in[761]
  PIN w_mask_in[762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.045 0.070 108.115 ;
    END
  END w_mask_in[762]
  PIN w_mask_in[763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.185 0.070 108.255 ;
    END
  END w_mask_in[763]
  PIN w_mask_in[764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END w_mask_in[764]
  PIN w_mask_in[765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.465 0.070 108.535 ;
    END
  END w_mask_in[765]
  PIN w_mask_in[766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.605 0.070 108.675 ;
    END
  END w_mask_in[766]
  PIN w_mask_in[767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END w_mask_in[767]
  PIN w_mask_in[768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.885 0.070 108.955 ;
    END
  END w_mask_in[768]
  PIN w_mask_in[769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.025 0.070 109.095 ;
    END
  END w_mask_in[769]
  PIN w_mask_in[770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END w_mask_in[770]
  PIN w_mask_in[771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.305 0.070 109.375 ;
    END
  END w_mask_in[771]
  PIN w_mask_in[772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.445 0.070 109.515 ;
    END
  END w_mask_in[772]
  PIN w_mask_in[773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.585 0.070 109.655 ;
    END
  END w_mask_in[773]
  PIN w_mask_in[774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.725 0.070 109.795 ;
    END
  END w_mask_in[774]
  PIN w_mask_in[775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.865 0.070 109.935 ;
    END
  END w_mask_in[775]
  PIN w_mask_in[776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.005 0.070 110.075 ;
    END
  END w_mask_in[776]
  PIN w_mask_in[777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.145 0.070 110.215 ;
    END
  END w_mask_in[777]
  PIN w_mask_in[778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.285 0.070 110.355 ;
    END
  END w_mask_in[778]
  PIN w_mask_in[779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.425 0.070 110.495 ;
    END
  END w_mask_in[779]
  PIN w_mask_in[780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.565 0.070 110.635 ;
    END
  END w_mask_in[780]
  PIN w_mask_in[781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.705 0.070 110.775 ;
    END
  END w_mask_in[781]
  PIN w_mask_in[782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END w_mask_in[782]
  PIN w_mask_in[783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.985 0.070 111.055 ;
    END
  END w_mask_in[783]
  PIN w_mask_in[784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.125 0.070 111.195 ;
    END
  END w_mask_in[784]
  PIN w_mask_in[785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.265 0.070 111.335 ;
    END
  END w_mask_in[785]
  PIN w_mask_in[786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.405 0.070 111.475 ;
    END
  END w_mask_in[786]
  PIN w_mask_in[787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.545 0.070 111.615 ;
    END
  END w_mask_in[787]
  PIN w_mask_in[788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.685 0.070 111.755 ;
    END
  END w_mask_in[788]
  PIN w_mask_in[789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.825 0.070 111.895 ;
    END
  END w_mask_in[789]
  PIN w_mask_in[790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.965 0.070 112.035 ;
    END
  END w_mask_in[790]
  PIN w_mask_in[791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.105 0.070 112.175 ;
    END
  END w_mask_in[791]
  PIN w_mask_in[792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END w_mask_in[792]
  PIN w_mask_in[793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.385 0.070 112.455 ;
    END
  END w_mask_in[793]
  PIN w_mask_in[794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.525 0.070 112.595 ;
    END
  END w_mask_in[794]
  PIN w_mask_in[795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.665 0.070 112.735 ;
    END
  END w_mask_in[795]
  PIN w_mask_in[796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.805 0.070 112.875 ;
    END
  END w_mask_in[796]
  PIN w_mask_in[797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.945 0.070 113.015 ;
    END
  END w_mask_in[797]
  PIN w_mask_in[798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END w_mask_in[798]
  PIN w_mask_in[799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.225 0.070 113.295 ;
    END
  END w_mask_in[799]
  PIN w_mask_in[800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.365 0.070 113.435 ;
    END
  END w_mask_in[800]
  PIN w_mask_in[801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.505 0.070 113.575 ;
    END
  END w_mask_in[801]
  PIN w_mask_in[802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.645 0.070 113.715 ;
    END
  END w_mask_in[802]
  PIN w_mask_in[803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.785 0.070 113.855 ;
    END
  END w_mask_in[803]
  PIN w_mask_in[804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.925 0.070 113.995 ;
    END
  END w_mask_in[804]
  PIN w_mask_in[805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.065 0.070 114.135 ;
    END
  END w_mask_in[805]
  PIN w_mask_in[806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.205 0.070 114.275 ;
    END
  END w_mask_in[806]
  PIN w_mask_in[807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.345 0.070 114.415 ;
    END
  END w_mask_in[807]
  PIN w_mask_in[808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.485 0.070 114.555 ;
    END
  END w_mask_in[808]
  PIN w_mask_in[809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.625 0.070 114.695 ;
    END
  END w_mask_in[809]
  PIN w_mask_in[810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.765 0.070 114.835 ;
    END
  END w_mask_in[810]
  PIN w_mask_in[811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.905 0.070 114.975 ;
    END
  END w_mask_in[811]
  PIN w_mask_in[812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END w_mask_in[812]
  PIN w_mask_in[813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.185 0.070 115.255 ;
    END
  END w_mask_in[813]
  PIN w_mask_in[814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END w_mask_in[814]
  PIN w_mask_in[815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.465 0.070 115.535 ;
    END
  END w_mask_in[815]
  PIN w_mask_in[816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.605 0.070 115.675 ;
    END
  END w_mask_in[816]
  PIN w_mask_in[817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.745 0.070 115.815 ;
    END
  END w_mask_in[817]
  PIN w_mask_in[818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.885 0.070 115.955 ;
    END
  END w_mask_in[818]
  PIN w_mask_in[819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.025 0.070 116.095 ;
    END
  END w_mask_in[819]
  PIN w_mask_in[820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END w_mask_in[820]
  PIN w_mask_in[821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.305 0.070 116.375 ;
    END
  END w_mask_in[821]
  PIN w_mask_in[822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.445 0.070 116.515 ;
    END
  END w_mask_in[822]
  PIN w_mask_in[823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.585 0.070 116.655 ;
    END
  END w_mask_in[823]
  PIN w_mask_in[824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.725 0.070 116.795 ;
    END
  END w_mask_in[824]
  PIN w_mask_in[825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.865 0.070 116.935 ;
    END
  END w_mask_in[825]
  PIN w_mask_in[826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END w_mask_in[826]
  PIN w_mask_in[827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.145 0.070 117.215 ;
    END
  END w_mask_in[827]
  PIN w_mask_in[828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.285 0.070 117.355 ;
    END
  END w_mask_in[828]
  PIN w_mask_in[829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.425 0.070 117.495 ;
    END
  END w_mask_in[829]
  PIN w_mask_in[830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END w_mask_in[830]
  PIN w_mask_in[831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.705 0.070 117.775 ;
    END
  END w_mask_in[831]
  PIN w_mask_in[832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.845 0.070 117.915 ;
    END
  END w_mask_in[832]
  PIN w_mask_in[833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.985 0.070 118.055 ;
    END
  END w_mask_in[833]
  PIN w_mask_in[834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END w_mask_in[834]
  PIN w_mask_in[835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.265 0.070 118.335 ;
    END
  END w_mask_in[835]
  PIN w_mask_in[836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.405 0.070 118.475 ;
    END
  END w_mask_in[836]
  PIN w_mask_in[837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.545 0.070 118.615 ;
    END
  END w_mask_in[837]
  PIN w_mask_in[838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.685 0.070 118.755 ;
    END
  END w_mask_in[838]
  PIN w_mask_in[839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.825 0.070 118.895 ;
    END
  END w_mask_in[839]
  PIN w_mask_in[840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END w_mask_in[840]
  PIN w_mask_in[841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.105 0.070 119.175 ;
    END
  END w_mask_in[841]
  PIN w_mask_in[842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.245 0.070 119.315 ;
    END
  END w_mask_in[842]
  PIN w_mask_in[843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.385 0.070 119.455 ;
    END
  END w_mask_in[843]
  PIN w_mask_in[844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.525 0.070 119.595 ;
    END
  END w_mask_in[844]
  PIN w_mask_in[845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.665 0.070 119.735 ;
    END
  END w_mask_in[845]
  PIN w_mask_in[846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END w_mask_in[846]
  PIN w_mask_in[847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.945 0.070 120.015 ;
    END
  END w_mask_in[847]
  PIN w_mask_in[848]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.085 0.070 120.155 ;
    END
  END w_mask_in[848]
  PIN w_mask_in[849]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.225 0.070 120.295 ;
    END
  END w_mask_in[849]
  PIN w_mask_in[850]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.365 0.070 120.435 ;
    END
  END w_mask_in[850]
  PIN w_mask_in[851]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.505 0.070 120.575 ;
    END
  END w_mask_in[851]
  PIN w_mask_in[852]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.645 0.070 120.715 ;
    END
  END w_mask_in[852]
  PIN w_mask_in[853]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.785 0.070 120.855 ;
    END
  END w_mask_in[853]
  PIN w_mask_in[854]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END w_mask_in[854]
  PIN w_mask_in[855]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.065 0.070 121.135 ;
    END
  END w_mask_in[855]
  PIN w_mask_in[856]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.205 0.070 121.275 ;
    END
  END w_mask_in[856]
  PIN w_mask_in[857]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.345 0.070 121.415 ;
    END
  END w_mask_in[857]
  PIN w_mask_in[858]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END w_mask_in[858]
  PIN w_mask_in[859]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.625 0.070 121.695 ;
    END
  END w_mask_in[859]
  PIN w_mask_in[860]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.765 0.070 121.835 ;
    END
  END w_mask_in[860]
  PIN w_mask_in[861]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.905 0.070 121.975 ;
    END
  END w_mask_in[861]
  PIN w_mask_in[862]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.045 0.070 122.115 ;
    END
  END w_mask_in[862]
  PIN w_mask_in[863]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.185 0.070 122.255 ;
    END
  END w_mask_in[863]
  PIN w_mask_in[864]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.325 0.070 122.395 ;
    END
  END w_mask_in[864]
  PIN w_mask_in[865]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.465 0.070 122.535 ;
    END
  END w_mask_in[865]
  PIN w_mask_in[866]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.605 0.070 122.675 ;
    END
  END w_mask_in[866]
  PIN w_mask_in[867]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.745 0.070 122.815 ;
    END
  END w_mask_in[867]
  PIN w_mask_in[868]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.885 0.070 122.955 ;
    END
  END w_mask_in[868]
  PIN w_mask_in[869]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.025 0.070 123.095 ;
    END
  END w_mask_in[869]
  PIN w_mask_in[870]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.165 0.070 123.235 ;
    END
  END w_mask_in[870]
  PIN w_mask_in[871]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.305 0.070 123.375 ;
    END
  END w_mask_in[871]
  PIN w_mask_in[872]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.445 0.070 123.515 ;
    END
  END w_mask_in[872]
  PIN w_mask_in[873]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.585 0.070 123.655 ;
    END
  END w_mask_in[873]
  PIN w_mask_in[874]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.725 0.070 123.795 ;
    END
  END w_mask_in[874]
  PIN w_mask_in[875]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.865 0.070 123.935 ;
    END
  END w_mask_in[875]
  PIN w_mask_in[876]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.005 0.070 124.075 ;
    END
  END w_mask_in[876]
  PIN w_mask_in[877]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.145 0.070 124.215 ;
    END
  END w_mask_in[877]
  PIN w_mask_in[878]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.285 0.070 124.355 ;
    END
  END w_mask_in[878]
  PIN w_mask_in[879]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.425 0.070 124.495 ;
    END
  END w_mask_in[879]
  PIN w_mask_in[880]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.565 0.070 124.635 ;
    END
  END w_mask_in[880]
  PIN w_mask_in[881]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.705 0.070 124.775 ;
    END
  END w_mask_in[881]
  PIN w_mask_in[882]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END w_mask_in[882]
  PIN w_mask_in[883]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.985 0.070 125.055 ;
    END
  END w_mask_in[883]
  PIN w_mask_in[884]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.125 0.070 125.195 ;
    END
  END w_mask_in[884]
  PIN w_mask_in[885]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.265 0.070 125.335 ;
    END
  END w_mask_in[885]
  PIN w_mask_in[886]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.405 0.070 125.475 ;
    END
  END w_mask_in[886]
  PIN w_mask_in[887]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.545 0.070 125.615 ;
    END
  END w_mask_in[887]
  PIN w_mask_in[888]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.685 0.070 125.755 ;
    END
  END w_mask_in[888]
  PIN w_mask_in[889]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.825 0.070 125.895 ;
    END
  END w_mask_in[889]
  PIN w_mask_in[890]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.965 0.070 126.035 ;
    END
  END w_mask_in[890]
  PIN w_mask_in[891]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.105 0.070 126.175 ;
    END
  END w_mask_in[891]
  PIN w_mask_in[892]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.245 0.070 126.315 ;
    END
  END w_mask_in[892]
  PIN w_mask_in[893]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.385 0.070 126.455 ;
    END
  END w_mask_in[893]
  PIN w_mask_in[894]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.525 0.070 126.595 ;
    END
  END w_mask_in[894]
  PIN w_mask_in[895]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.665 0.070 126.735 ;
    END
  END w_mask_in[895]
  PIN w_mask_in[896]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.805 0.070 126.875 ;
    END
  END w_mask_in[896]
  PIN w_mask_in[897]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.945 0.070 127.015 ;
    END
  END w_mask_in[897]
  PIN w_mask_in[898]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.085 0.070 127.155 ;
    END
  END w_mask_in[898]
  PIN w_mask_in[899]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.225 0.070 127.295 ;
    END
  END w_mask_in[899]
  PIN w_mask_in[900]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.365 0.070 127.435 ;
    END
  END w_mask_in[900]
  PIN w_mask_in[901]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.505 0.070 127.575 ;
    END
  END w_mask_in[901]
  PIN w_mask_in[902]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.645 0.070 127.715 ;
    END
  END w_mask_in[902]
  PIN w_mask_in[903]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.785 0.070 127.855 ;
    END
  END w_mask_in[903]
  PIN w_mask_in[904]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.925 0.070 127.995 ;
    END
  END w_mask_in[904]
  PIN w_mask_in[905]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.065 0.070 128.135 ;
    END
  END w_mask_in[905]
  PIN w_mask_in[906]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.205 0.070 128.275 ;
    END
  END w_mask_in[906]
  PIN w_mask_in[907]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.345 0.070 128.415 ;
    END
  END w_mask_in[907]
  PIN w_mask_in[908]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.485 0.070 128.555 ;
    END
  END w_mask_in[908]
  PIN w_mask_in[909]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.625 0.070 128.695 ;
    END
  END w_mask_in[909]
  PIN w_mask_in[910]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END w_mask_in[910]
  PIN w_mask_in[911]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.905 0.070 128.975 ;
    END
  END w_mask_in[911]
  PIN w_mask_in[912]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.045 0.070 129.115 ;
    END
  END w_mask_in[912]
  PIN w_mask_in[913]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.185 0.070 129.255 ;
    END
  END w_mask_in[913]
  PIN w_mask_in[914]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END w_mask_in[914]
  PIN w_mask_in[915]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.465 0.070 129.535 ;
    END
  END w_mask_in[915]
  PIN w_mask_in[916]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.605 0.070 129.675 ;
    END
  END w_mask_in[916]
  PIN w_mask_in[917]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.745 0.070 129.815 ;
    END
  END w_mask_in[917]
  PIN w_mask_in[918]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END w_mask_in[918]
  PIN w_mask_in[919]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.025 0.070 130.095 ;
    END
  END w_mask_in[919]
  PIN w_mask_in[920]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.165 0.070 130.235 ;
    END
  END w_mask_in[920]
  PIN w_mask_in[921]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.305 0.070 130.375 ;
    END
  END w_mask_in[921]
  PIN w_mask_in[922]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.445 0.070 130.515 ;
    END
  END w_mask_in[922]
  PIN w_mask_in[923]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.585 0.070 130.655 ;
    END
  END w_mask_in[923]
  PIN w_mask_in[924]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END w_mask_in[924]
  PIN w_mask_in[925]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.865 0.070 130.935 ;
    END
  END w_mask_in[925]
  PIN w_mask_in[926]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.005 0.070 131.075 ;
    END
  END w_mask_in[926]
  PIN w_mask_in[927]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.145 0.070 131.215 ;
    END
  END w_mask_in[927]
  PIN w_mask_in[928]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.285 0.070 131.355 ;
    END
  END w_mask_in[928]
  PIN w_mask_in[929]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.425 0.070 131.495 ;
    END
  END w_mask_in[929]
  PIN w_mask_in[930]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.565 0.070 131.635 ;
    END
  END w_mask_in[930]
  PIN w_mask_in[931]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.705 0.070 131.775 ;
    END
  END w_mask_in[931]
  PIN w_mask_in[932]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.845 0.070 131.915 ;
    END
  END w_mask_in[932]
  PIN w_mask_in[933]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.985 0.070 132.055 ;
    END
  END w_mask_in[933]
  PIN w_mask_in[934]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.125 0.070 132.195 ;
    END
  END w_mask_in[934]
  PIN w_mask_in[935]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.265 0.070 132.335 ;
    END
  END w_mask_in[935]
  PIN w_mask_in[936]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.405 0.070 132.475 ;
    END
  END w_mask_in[936]
  PIN w_mask_in[937]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.545 0.070 132.615 ;
    END
  END w_mask_in[937]
  PIN w_mask_in[938]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.685 0.070 132.755 ;
    END
  END w_mask_in[938]
  PIN w_mask_in[939]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.825 0.070 132.895 ;
    END
  END w_mask_in[939]
  PIN w_mask_in[940]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.965 0.070 133.035 ;
    END
  END w_mask_in[940]
  PIN w_mask_in[941]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.105 0.070 133.175 ;
    END
  END w_mask_in[941]
  PIN w_mask_in[942]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.245 0.070 133.315 ;
    END
  END w_mask_in[942]
  PIN w_mask_in[943]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.385 0.070 133.455 ;
    END
  END w_mask_in[943]
  PIN w_mask_in[944]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.525 0.070 133.595 ;
    END
  END w_mask_in[944]
  PIN w_mask_in[945]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.665 0.070 133.735 ;
    END
  END w_mask_in[945]
  PIN w_mask_in[946]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.805 0.070 133.875 ;
    END
  END w_mask_in[946]
  PIN w_mask_in[947]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.945 0.070 134.015 ;
    END
  END w_mask_in[947]
  PIN w_mask_in[948]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.085 0.070 134.155 ;
    END
  END w_mask_in[948]
  PIN w_mask_in[949]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.225 0.070 134.295 ;
    END
  END w_mask_in[949]
  PIN w_mask_in[950]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.365 0.070 134.435 ;
    END
  END w_mask_in[950]
  PIN w_mask_in[951]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.505 0.070 134.575 ;
    END
  END w_mask_in[951]
  PIN w_mask_in[952]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.645 0.070 134.715 ;
    END
  END w_mask_in[952]
  PIN w_mask_in[953]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.785 0.070 134.855 ;
    END
  END w_mask_in[953]
  PIN w_mask_in[954]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END w_mask_in[954]
  PIN w_mask_in[955]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.065 0.070 135.135 ;
    END
  END w_mask_in[955]
  PIN w_mask_in[956]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.205 0.070 135.275 ;
    END
  END w_mask_in[956]
  PIN w_mask_in[957]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.345 0.070 135.415 ;
    END
  END w_mask_in[957]
  PIN w_mask_in[958]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.485 0.070 135.555 ;
    END
  END w_mask_in[958]
  PIN w_mask_in[959]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.625 0.070 135.695 ;
    END
  END w_mask_in[959]
  PIN w_mask_in[960]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.765 0.070 135.835 ;
    END
  END w_mask_in[960]
  PIN w_mask_in[961]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.905 0.070 135.975 ;
    END
  END w_mask_in[961]
  PIN w_mask_in[962]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.045 0.070 136.115 ;
    END
  END w_mask_in[962]
  PIN w_mask_in[963]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.185 0.070 136.255 ;
    END
  END w_mask_in[963]
  PIN w_mask_in[964]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.325 0.070 136.395 ;
    END
  END w_mask_in[964]
  PIN w_mask_in[965]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.465 0.070 136.535 ;
    END
  END w_mask_in[965]
  PIN w_mask_in[966]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END w_mask_in[966]
  PIN w_mask_in[967]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.745 0.070 136.815 ;
    END
  END w_mask_in[967]
  PIN w_mask_in[968]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.885 0.070 136.955 ;
    END
  END w_mask_in[968]
  PIN w_mask_in[969]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.025 0.070 137.095 ;
    END
  END w_mask_in[969]
  PIN w_mask_in[970]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.165 0.070 137.235 ;
    END
  END w_mask_in[970]
  PIN w_mask_in[971]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.305 0.070 137.375 ;
    END
  END w_mask_in[971]
  PIN w_mask_in[972]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.445 0.070 137.515 ;
    END
  END w_mask_in[972]
  PIN w_mask_in[973]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.585 0.070 137.655 ;
    END
  END w_mask_in[973]
  PIN w_mask_in[974]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.725 0.070 137.795 ;
    END
  END w_mask_in[974]
  PIN w_mask_in[975]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.865 0.070 137.935 ;
    END
  END w_mask_in[975]
  PIN w_mask_in[976]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.005 0.070 138.075 ;
    END
  END w_mask_in[976]
  PIN w_mask_in[977]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.145 0.070 138.215 ;
    END
  END w_mask_in[977]
  PIN w_mask_in[978]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END w_mask_in[978]
  PIN w_mask_in[979]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.425 0.070 138.495 ;
    END
  END w_mask_in[979]
  PIN w_mask_in[980]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.565 0.070 138.635 ;
    END
  END w_mask_in[980]
  PIN w_mask_in[981]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.705 0.070 138.775 ;
    END
  END w_mask_in[981]
  PIN w_mask_in[982]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.845 0.070 138.915 ;
    END
  END w_mask_in[982]
  PIN w_mask_in[983]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.985 0.070 139.055 ;
    END
  END w_mask_in[983]
  PIN w_mask_in[984]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END w_mask_in[984]
  PIN w_mask_in[985]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.265 0.070 139.335 ;
    END
  END w_mask_in[985]
  PIN w_mask_in[986]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.405 0.070 139.475 ;
    END
  END w_mask_in[986]
  PIN w_mask_in[987]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.545 0.070 139.615 ;
    END
  END w_mask_in[987]
  PIN w_mask_in[988]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.685 0.070 139.755 ;
    END
  END w_mask_in[988]
  PIN w_mask_in[989]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.825 0.070 139.895 ;
    END
  END w_mask_in[989]
  PIN w_mask_in[990]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END w_mask_in[990]
  PIN w_mask_in[991]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.105 0.070 140.175 ;
    END
  END w_mask_in[991]
  PIN w_mask_in[992]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.245 0.070 140.315 ;
    END
  END w_mask_in[992]
  PIN w_mask_in[993]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.385 0.070 140.455 ;
    END
  END w_mask_in[993]
  PIN w_mask_in[994]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.525 0.070 140.595 ;
    END
  END w_mask_in[994]
  PIN w_mask_in[995]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.665 0.070 140.735 ;
    END
  END w_mask_in[995]
  PIN w_mask_in[996]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.805 0.070 140.875 ;
    END
  END w_mask_in[996]
  PIN w_mask_in[997]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.945 0.070 141.015 ;
    END
  END w_mask_in[997]
  PIN w_mask_in[998]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.085 0.070 141.155 ;
    END
  END w_mask_in[998]
  PIN w_mask_in[999]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.225 0.070 141.295 ;
    END
  END w_mask_in[999]
  PIN w_mask_in[1000]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.365 0.070 141.435 ;
    END
  END w_mask_in[1000]
  PIN w_mask_in[1001]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.505 0.070 141.575 ;
    END
  END w_mask_in[1001]
  PIN w_mask_in[1002]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END w_mask_in[1002]
  PIN w_mask_in[1003]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.785 0.070 141.855 ;
    END
  END w_mask_in[1003]
  PIN w_mask_in[1004]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.925 0.070 141.995 ;
    END
  END w_mask_in[1004]
  PIN w_mask_in[1005]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.065 0.070 142.135 ;
    END
  END w_mask_in[1005]
  PIN w_mask_in[1006]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.205 0.070 142.275 ;
    END
  END w_mask_in[1006]
  PIN w_mask_in[1007]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.345 0.070 142.415 ;
    END
  END w_mask_in[1007]
  PIN w_mask_in[1008]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END w_mask_in[1008]
  PIN w_mask_in[1009]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.625 0.070 142.695 ;
    END
  END w_mask_in[1009]
  PIN w_mask_in[1010]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.765 0.070 142.835 ;
    END
  END w_mask_in[1010]
  PIN w_mask_in[1011]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.905 0.070 142.975 ;
    END
  END w_mask_in[1011]
  PIN w_mask_in[1012]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.045 0.070 143.115 ;
    END
  END w_mask_in[1012]
  PIN w_mask_in[1013]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.185 0.070 143.255 ;
    END
  END w_mask_in[1013]
  PIN w_mask_in[1014]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END w_mask_in[1014]
  PIN w_mask_in[1015]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.465 0.070 143.535 ;
    END
  END w_mask_in[1015]
  PIN w_mask_in[1016]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.605 0.070 143.675 ;
    END
  END w_mask_in[1016]
  PIN w_mask_in[1017]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.745 0.070 143.815 ;
    END
  END w_mask_in[1017]
  PIN w_mask_in[1018]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.885 0.070 143.955 ;
    END
  END w_mask_in[1018]
  PIN w_mask_in[1019]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.025 0.070 144.095 ;
    END
  END w_mask_in[1019]
  PIN w_mask_in[1020]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.165 0.070 144.235 ;
    END
  END w_mask_in[1020]
  PIN w_mask_in[1021]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.305 0.070 144.375 ;
    END
  END w_mask_in[1021]
  PIN w_mask_in[1022]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END w_mask_in[1022]
  PIN w_mask_in[1023]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.585 0.070 144.655 ;
    END
  END w_mask_in[1023]
  PIN w_mask_in[1024]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.725 0.070 144.795 ;
    END
  END w_mask_in[1024]
  PIN w_mask_in[1025]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.865 0.070 144.935 ;
    END
  END w_mask_in[1025]
  PIN w_mask_in[1026]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END w_mask_in[1026]
  PIN w_mask_in[1027]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.145 0.070 145.215 ;
    END
  END w_mask_in[1027]
  PIN w_mask_in[1028]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.285 0.070 145.355 ;
    END
  END w_mask_in[1028]
  PIN w_mask_in[1029]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.425 0.070 145.495 ;
    END
  END w_mask_in[1029]
  PIN w_mask_in[1030]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.565 0.070 145.635 ;
    END
  END w_mask_in[1030]
  PIN w_mask_in[1031]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.705 0.070 145.775 ;
    END
  END w_mask_in[1031]
  PIN w_mask_in[1032]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.845 0.070 145.915 ;
    END
  END w_mask_in[1032]
  PIN w_mask_in[1033]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.985 0.070 146.055 ;
    END
  END w_mask_in[1033]
  PIN w_mask_in[1034]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.125 0.070 146.195 ;
    END
  END w_mask_in[1034]
  PIN w_mask_in[1035]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.265 0.070 146.335 ;
    END
  END w_mask_in[1035]
  PIN w_mask_in[1036]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.405 0.070 146.475 ;
    END
  END w_mask_in[1036]
  PIN w_mask_in[1037]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.545 0.070 146.615 ;
    END
  END w_mask_in[1037]
  PIN w_mask_in[1038]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END w_mask_in[1038]
  PIN w_mask_in[1039]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.825 0.070 146.895 ;
    END
  END w_mask_in[1039]
  PIN w_mask_in[1040]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.965 0.070 147.035 ;
    END
  END w_mask_in[1040]
  PIN w_mask_in[1041]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.105 0.070 147.175 ;
    END
  END w_mask_in[1041]
  PIN w_mask_in[1042]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.245 0.070 147.315 ;
    END
  END w_mask_in[1042]
  PIN w_mask_in[1043]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.385 0.070 147.455 ;
    END
  END w_mask_in[1043]
  PIN w_mask_in[1044]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.525 0.070 147.595 ;
    END
  END w_mask_in[1044]
  PIN w_mask_in[1045]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.665 0.070 147.735 ;
    END
  END w_mask_in[1045]
  PIN w_mask_in[1046]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.805 0.070 147.875 ;
    END
  END w_mask_in[1046]
  PIN w_mask_in[1047]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.945 0.070 148.015 ;
    END
  END w_mask_in[1047]
  PIN w_mask_in[1048]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.085 0.070 148.155 ;
    END
  END w_mask_in[1048]
  PIN w_mask_in[1049]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.225 0.070 148.295 ;
    END
  END w_mask_in[1049]
  PIN w_mask_in[1050]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END w_mask_in[1050]
  PIN w_mask_in[1051]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.505 0.070 148.575 ;
    END
  END w_mask_in[1051]
  PIN w_mask_in[1052]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.645 0.070 148.715 ;
    END
  END w_mask_in[1052]
  PIN w_mask_in[1053]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.785 0.070 148.855 ;
    END
  END w_mask_in[1053]
  PIN w_mask_in[1054]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.925 0.070 148.995 ;
    END
  END w_mask_in[1054]
  PIN w_mask_in[1055]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.065 0.070 149.135 ;
    END
  END w_mask_in[1055]
  PIN w_mask_in[1056]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.205 0.070 149.275 ;
    END
  END w_mask_in[1056]
  PIN w_mask_in[1057]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.345 0.070 149.415 ;
    END
  END w_mask_in[1057]
  PIN w_mask_in[1058]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.485 0.070 149.555 ;
    END
  END w_mask_in[1058]
  PIN w_mask_in[1059]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.625 0.070 149.695 ;
    END
  END w_mask_in[1059]
  PIN w_mask_in[1060]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.765 0.070 149.835 ;
    END
  END w_mask_in[1060]
  PIN w_mask_in[1061]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.905 0.070 149.975 ;
    END
  END w_mask_in[1061]
  PIN w_mask_in[1062]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.045 0.070 150.115 ;
    END
  END w_mask_in[1062]
  PIN w_mask_in[1063]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.185 0.070 150.255 ;
    END
  END w_mask_in[1063]
  PIN w_mask_in[1064]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END w_mask_in[1064]
  PIN w_mask_in[1065]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.465 0.070 150.535 ;
    END
  END w_mask_in[1065]
  PIN w_mask_in[1066]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END w_mask_in[1066]
  PIN w_mask_in[1067]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.745 0.070 150.815 ;
    END
  END w_mask_in[1067]
  PIN w_mask_in[1068]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.885 0.070 150.955 ;
    END
  END w_mask_in[1068]
  PIN w_mask_in[1069]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.025 0.070 151.095 ;
    END
  END w_mask_in[1069]
  PIN w_mask_in[1070]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.165 0.070 151.235 ;
    END
  END w_mask_in[1070]
  PIN w_mask_in[1071]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.305 0.070 151.375 ;
    END
  END w_mask_in[1071]
  PIN w_mask_in[1072]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.445 0.070 151.515 ;
    END
  END w_mask_in[1072]
  PIN w_mask_in[1073]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.585 0.070 151.655 ;
    END
  END w_mask_in[1073]
  PIN w_mask_in[1074]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.725 0.070 151.795 ;
    END
  END w_mask_in[1074]
  PIN w_mask_in[1075]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.865 0.070 151.935 ;
    END
  END w_mask_in[1075]
  PIN w_mask_in[1076]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.005 0.070 152.075 ;
    END
  END w_mask_in[1076]
  PIN w_mask_in[1077]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.145 0.070 152.215 ;
    END
  END w_mask_in[1077]
  PIN w_mask_in[1078]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END w_mask_in[1078]
  PIN w_mask_in[1079]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.425 0.070 152.495 ;
    END
  END w_mask_in[1079]
  PIN w_mask_in[1080]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.565 0.070 152.635 ;
    END
  END w_mask_in[1080]
  PIN w_mask_in[1081]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.705 0.070 152.775 ;
    END
  END w_mask_in[1081]
  PIN w_mask_in[1082]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.845 0.070 152.915 ;
    END
  END w_mask_in[1082]
  PIN w_mask_in[1083]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.985 0.070 153.055 ;
    END
  END w_mask_in[1083]
  PIN w_mask_in[1084]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.125 0.070 153.195 ;
    END
  END w_mask_in[1084]
  PIN w_mask_in[1085]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.265 0.070 153.335 ;
    END
  END w_mask_in[1085]
  PIN w_mask_in[1086]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.405 0.070 153.475 ;
    END
  END w_mask_in[1086]
  PIN w_mask_in[1087]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.545 0.070 153.615 ;
    END
  END w_mask_in[1087]
  PIN w_mask_in[1088]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.685 0.070 153.755 ;
    END
  END w_mask_in[1088]
  PIN w_mask_in[1089]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.825 0.070 153.895 ;
    END
  END w_mask_in[1089]
  PIN w_mask_in[1090]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.965 0.070 154.035 ;
    END
  END w_mask_in[1090]
  PIN w_mask_in[1091]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.105 0.070 154.175 ;
    END
  END w_mask_in[1091]
  PIN w_mask_in[1092]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END w_mask_in[1092]
  PIN w_mask_in[1093]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.385 0.070 154.455 ;
    END
  END w_mask_in[1093]
  PIN w_mask_in[1094]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END w_mask_in[1094]
  PIN w_mask_in[1095]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.665 0.070 154.735 ;
    END
  END w_mask_in[1095]
  PIN w_mask_in[1096]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.805 0.070 154.875 ;
    END
  END w_mask_in[1096]
  PIN w_mask_in[1097]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.945 0.070 155.015 ;
    END
  END w_mask_in[1097]
  PIN w_mask_in[1098]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.085 0.070 155.155 ;
    END
  END w_mask_in[1098]
  PIN w_mask_in[1099]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.225 0.070 155.295 ;
    END
  END w_mask_in[1099]
  PIN w_mask_in[1100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.365 0.070 155.435 ;
    END
  END w_mask_in[1100]
  PIN w_mask_in[1101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.505 0.070 155.575 ;
    END
  END w_mask_in[1101]
  PIN w_mask_in[1102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.645 0.070 155.715 ;
    END
  END w_mask_in[1102]
  PIN w_mask_in[1103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.785 0.070 155.855 ;
    END
  END w_mask_in[1103]
  PIN w_mask_in[1104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.925 0.070 155.995 ;
    END
  END w_mask_in[1104]
  PIN w_mask_in[1105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.065 0.070 156.135 ;
    END
  END w_mask_in[1105]
  PIN w_mask_in[1106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.205 0.070 156.275 ;
    END
  END w_mask_in[1106]
  PIN w_mask_in[1107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.345 0.070 156.415 ;
    END
  END w_mask_in[1107]
  PIN w_mask_in[1108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.485 0.070 156.555 ;
    END
  END w_mask_in[1108]
  PIN w_mask_in[1109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.625 0.070 156.695 ;
    END
  END w_mask_in[1109]
  PIN w_mask_in[1110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.765 0.070 156.835 ;
    END
  END w_mask_in[1110]
  PIN w_mask_in[1111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.905 0.070 156.975 ;
    END
  END w_mask_in[1111]
  PIN w_mask_in[1112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.045 0.070 157.115 ;
    END
  END w_mask_in[1112]
  PIN w_mask_in[1113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.185 0.070 157.255 ;
    END
  END w_mask_in[1113]
  PIN w_mask_in[1114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.325 0.070 157.395 ;
    END
  END w_mask_in[1114]
  PIN w_mask_in[1115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.465 0.070 157.535 ;
    END
  END w_mask_in[1115]
  PIN w_mask_in[1116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.605 0.070 157.675 ;
    END
  END w_mask_in[1116]
  PIN w_mask_in[1117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.745 0.070 157.815 ;
    END
  END w_mask_in[1117]
  PIN w_mask_in[1118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.885 0.070 157.955 ;
    END
  END w_mask_in[1118]
  PIN w_mask_in[1119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.025 0.070 158.095 ;
    END
  END w_mask_in[1119]
  PIN w_mask_in[1120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.165 0.070 158.235 ;
    END
  END w_mask_in[1120]
  PIN w_mask_in[1121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.305 0.070 158.375 ;
    END
  END w_mask_in[1121]
  PIN w_mask_in[1122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.445 0.070 158.515 ;
    END
  END w_mask_in[1122]
  PIN w_mask_in[1123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.585 0.070 158.655 ;
    END
  END w_mask_in[1123]
  PIN w_mask_in[1124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.725 0.070 158.795 ;
    END
  END w_mask_in[1124]
  PIN w_mask_in[1125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.865 0.070 158.935 ;
    END
  END w_mask_in[1125]
  PIN w_mask_in[1126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.005 0.070 159.075 ;
    END
  END w_mask_in[1126]
  PIN w_mask_in[1127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.145 0.070 159.215 ;
    END
  END w_mask_in[1127]
  PIN w_mask_in[1128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.285 0.070 159.355 ;
    END
  END w_mask_in[1128]
  PIN w_mask_in[1129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.425 0.070 159.495 ;
    END
  END w_mask_in[1129]
  PIN w_mask_in[1130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.565 0.070 159.635 ;
    END
  END w_mask_in[1130]
  PIN w_mask_in[1131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.705 0.070 159.775 ;
    END
  END w_mask_in[1131]
  PIN w_mask_in[1132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.845 0.070 159.915 ;
    END
  END w_mask_in[1132]
  PIN w_mask_in[1133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.985 0.070 160.055 ;
    END
  END w_mask_in[1133]
  PIN w_mask_in[1134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END w_mask_in[1134]
  PIN w_mask_in[1135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.265 0.070 160.335 ;
    END
  END w_mask_in[1135]
  PIN w_mask_in[1136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.405 0.070 160.475 ;
    END
  END w_mask_in[1136]
  PIN w_mask_in[1137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.545 0.070 160.615 ;
    END
  END w_mask_in[1137]
  PIN w_mask_in[1138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.685 0.070 160.755 ;
    END
  END w_mask_in[1138]
  PIN w_mask_in[1139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.825 0.070 160.895 ;
    END
  END w_mask_in[1139]
  PIN w_mask_in[1140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.965 0.070 161.035 ;
    END
  END w_mask_in[1140]
  PIN w_mask_in[1141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.105 0.070 161.175 ;
    END
  END w_mask_in[1141]
  PIN w_mask_in[1142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.245 0.070 161.315 ;
    END
  END w_mask_in[1142]
  PIN w_mask_in[1143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.385 0.070 161.455 ;
    END
  END w_mask_in[1143]
  PIN w_mask_in[1144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.525 0.070 161.595 ;
    END
  END w_mask_in[1144]
  PIN w_mask_in[1145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.665 0.070 161.735 ;
    END
  END w_mask_in[1145]
  PIN w_mask_in[1146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.805 0.070 161.875 ;
    END
  END w_mask_in[1146]
  PIN w_mask_in[1147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.945 0.070 162.015 ;
    END
  END w_mask_in[1147]
  PIN w_mask_in[1148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.085 0.070 162.155 ;
    END
  END w_mask_in[1148]
  PIN w_mask_in[1149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.225 0.070 162.295 ;
    END
  END w_mask_in[1149]
  PIN w_mask_in[1150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.365 0.070 162.435 ;
    END
  END w_mask_in[1150]
  PIN w_mask_in[1151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.505 0.070 162.575 ;
    END
  END w_mask_in[1151]
  PIN w_mask_in[1152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.645 0.070 162.715 ;
    END
  END w_mask_in[1152]
  PIN w_mask_in[1153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.785 0.070 162.855 ;
    END
  END w_mask_in[1153]
  PIN w_mask_in[1154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.925 0.070 162.995 ;
    END
  END w_mask_in[1154]
  PIN w_mask_in[1155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.065 0.070 163.135 ;
    END
  END w_mask_in[1155]
  PIN w_mask_in[1156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.205 0.070 163.275 ;
    END
  END w_mask_in[1156]
  PIN w_mask_in[1157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.345 0.070 163.415 ;
    END
  END w_mask_in[1157]
  PIN w_mask_in[1158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.485 0.070 163.555 ;
    END
  END w_mask_in[1158]
  PIN w_mask_in[1159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.625 0.070 163.695 ;
    END
  END w_mask_in[1159]
  PIN w_mask_in[1160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.765 0.070 163.835 ;
    END
  END w_mask_in[1160]
  PIN w_mask_in[1161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.905 0.070 163.975 ;
    END
  END w_mask_in[1161]
  PIN w_mask_in[1162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.045 0.070 164.115 ;
    END
  END w_mask_in[1162]
  PIN w_mask_in[1163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.185 0.070 164.255 ;
    END
  END w_mask_in[1163]
  PIN w_mask_in[1164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.325 0.070 164.395 ;
    END
  END w_mask_in[1164]
  PIN w_mask_in[1165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.465 0.070 164.535 ;
    END
  END w_mask_in[1165]
  PIN w_mask_in[1166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.605 0.070 164.675 ;
    END
  END w_mask_in[1166]
  PIN w_mask_in[1167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.745 0.070 164.815 ;
    END
  END w_mask_in[1167]
  PIN w_mask_in[1168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.885 0.070 164.955 ;
    END
  END w_mask_in[1168]
  PIN w_mask_in[1169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.025 0.070 165.095 ;
    END
  END w_mask_in[1169]
  PIN w_mask_in[1170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END w_mask_in[1170]
  PIN w_mask_in[1171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.305 0.070 165.375 ;
    END
  END w_mask_in[1171]
  PIN w_mask_in[1172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.445 0.070 165.515 ;
    END
  END w_mask_in[1172]
  PIN w_mask_in[1173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.585 0.070 165.655 ;
    END
  END w_mask_in[1173]
  PIN w_mask_in[1174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.725 0.070 165.795 ;
    END
  END w_mask_in[1174]
  PIN w_mask_in[1175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.865 0.070 165.935 ;
    END
  END w_mask_in[1175]
  PIN w_mask_in[1176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.005 0.070 166.075 ;
    END
  END w_mask_in[1176]
  PIN w_mask_in[1177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.145 0.070 166.215 ;
    END
  END w_mask_in[1177]
  PIN w_mask_in[1178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.285 0.070 166.355 ;
    END
  END w_mask_in[1178]
  PIN w_mask_in[1179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.425 0.070 166.495 ;
    END
  END w_mask_in[1179]
  PIN w_mask_in[1180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.565 0.070 166.635 ;
    END
  END w_mask_in[1180]
  PIN w_mask_in[1181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.705 0.070 166.775 ;
    END
  END w_mask_in[1181]
  PIN w_mask_in[1182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.845 0.070 166.915 ;
    END
  END w_mask_in[1182]
  PIN w_mask_in[1183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.985 0.070 167.055 ;
    END
  END w_mask_in[1183]
  PIN w_mask_in[1184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.125 0.070 167.195 ;
    END
  END w_mask_in[1184]
  PIN w_mask_in[1185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.265 0.070 167.335 ;
    END
  END w_mask_in[1185]
  PIN w_mask_in[1186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.405 0.070 167.475 ;
    END
  END w_mask_in[1186]
  PIN w_mask_in[1187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.545 0.070 167.615 ;
    END
  END w_mask_in[1187]
  PIN w_mask_in[1188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END w_mask_in[1188]
  PIN w_mask_in[1189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.825 0.070 167.895 ;
    END
  END w_mask_in[1189]
  PIN w_mask_in[1190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.965 0.070 168.035 ;
    END
  END w_mask_in[1190]
  PIN w_mask_in[1191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.105 0.070 168.175 ;
    END
  END w_mask_in[1191]
  PIN w_mask_in[1192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.245 0.070 168.315 ;
    END
  END w_mask_in[1192]
  PIN w_mask_in[1193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.385 0.070 168.455 ;
    END
  END w_mask_in[1193]
  PIN w_mask_in[1194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.525 0.070 168.595 ;
    END
  END w_mask_in[1194]
  PIN w_mask_in[1195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.665 0.070 168.735 ;
    END
  END w_mask_in[1195]
  PIN w_mask_in[1196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.805 0.070 168.875 ;
    END
  END w_mask_in[1196]
  PIN w_mask_in[1197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.945 0.070 169.015 ;
    END
  END w_mask_in[1197]
  PIN w_mask_in[1198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.085 0.070 169.155 ;
    END
  END w_mask_in[1198]
  PIN w_mask_in[1199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.225 0.070 169.295 ;
    END
  END w_mask_in[1199]
  PIN w_mask_in[1200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.365 0.070 169.435 ;
    END
  END w_mask_in[1200]
  PIN w_mask_in[1201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.505 0.070 169.575 ;
    END
  END w_mask_in[1201]
  PIN w_mask_in[1202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.645 0.070 169.715 ;
    END
  END w_mask_in[1202]
  PIN w_mask_in[1203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.785 0.070 169.855 ;
    END
  END w_mask_in[1203]
  PIN w_mask_in[1204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.925 0.070 169.995 ;
    END
  END w_mask_in[1204]
  PIN w_mask_in[1205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.065 0.070 170.135 ;
    END
  END w_mask_in[1205]
  PIN w_mask_in[1206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END w_mask_in[1206]
  PIN w_mask_in[1207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.345 0.070 170.415 ;
    END
  END w_mask_in[1207]
  PIN w_mask_in[1208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.485 0.070 170.555 ;
    END
  END w_mask_in[1208]
  PIN w_mask_in[1209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.625 0.070 170.695 ;
    END
  END w_mask_in[1209]
  PIN w_mask_in[1210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.765 0.070 170.835 ;
    END
  END w_mask_in[1210]
  PIN w_mask_in[1211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.905 0.070 170.975 ;
    END
  END w_mask_in[1211]
  PIN w_mask_in[1212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.045 0.070 171.115 ;
    END
  END w_mask_in[1212]
  PIN w_mask_in[1213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.185 0.070 171.255 ;
    END
  END w_mask_in[1213]
  PIN w_mask_in[1214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.325 0.070 171.395 ;
    END
  END w_mask_in[1214]
  PIN w_mask_in[1215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.465 0.070 171.535 ;
    END
  END w_mask_in[1215]
  PIN w_mask_in[1216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.605 0.070 171.675 ;
    END
  END w_mask_in[1216]
  PIN w_mask_in[1217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.745 0.070 171.815 ;
    END
  END w_mask_in[1217]
  PIN w_mask_in[1218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END w_mask_in[1218]
  PIN w_mask_in[1219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.025 0.070 172.095 ;
    END
  END w_mask_in[1219]
  PIN w_mask_in[1220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END w_mask_in[1220]
  PIN w_mask_in[1221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.305 0.070 172.375 ;
    END
  END w_mask_in[1221]
  PIN w_mask_in[1222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.445 0.070 172.515 ;
    END
  END w_mask_in[1222]
  PIN w_mask_in[1223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.585 0.070 172.655 ;
    END
  END w_mask_in[1223]
  PIN w_mask_in[1224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.725 0.070 172.795 ;
    END
  END w_mask_in[1224]
  PIN w_mask_in[1225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.865 0.070 172.935 ;
    END
  END w_mask_in[1225]
  PIN w_mask_in[1226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.005 0.070 173.075 ;
    END
  END w_mask_in[1226]
  PIN w_mask_in[1227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.145 0.070 173.215 ;
    END
  END w_mask_in[1227]
  PIN w_mask_in[1228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.285 0.070 173.355 ;
    END
  END w_mask_in[1228]
  PIN w_mask_in[1229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.425 0.070 173.495 ;
    END
  END w_mask_in[1229]
  PIN w_mask_in[1230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.565 0.070 173.635 ;
    END
  END w_mask_in[1230]
  PIN w_mask_in[1231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.705 0.070 173.775 ;
    END
  END w_mask_in[1231]
  PIN w_mask_in[1232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.845 0.070 173.915 ;
    END
  END w_mask_in[1232]
  PIN w_mask_in[1233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.985 0.070 174.055 ;
    END
  END w_mask_in[1233]
  PIN w_mask_in[1234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.125 0.070 174.195 ;
    END
  END w_mask_in[1234]
  PIN w_mask_in[1235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.265 0.070 174.335 ;
    END
  END w_mask_in[1235]
  PIN w_mask_in[1236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.405 0.070 174.475 ;
    END
  END w_mask_in[1236]
  PIN w_mask_in[1237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.545 0.070 174.615 ;
    END
  END w_mask_in[1237]
  PIN w_mask_in[1238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.685 0.070 174.755 ;
    END
  END w_mask_in[1238]
  PIN w_mask_in[1239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.825 0.070 174.895 ;
    END
  END w_mask_in[1239]
  PIN w_mask_in[1240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.965 0.070 175.035 ;
    END
  END w_mask_in[1240]
  PIN w_mask_in[1241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.105 0.070 175.175 ;
    END
  END w_mask_in[1241]
  PIN w_mask_in[1242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.245 0.070 175.315 ;
    END
  END w_mask_in[1242]
  PIN w_mask_in[1243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.385 0.070 175.455 ;
    END
  END w_mask_in[1243]
  PIN w_mask_in[1244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.525 0.070 175.595 ;
    END
  END w_mask_in[1244]
  PIN w_mask_in[1245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.665 0.070 175.735 ;
    END
  END w_mask_in[1245]
  PIN w_mask_in[1246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.805 0.070 175.875 ;
    END
  END w_mask_in[1246]
  PIN w_mask_in[1247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.945 0.070 176.015 ;
    END
  END w_mask_in[1247]
  PIN w_mask_in[1248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.085 0.070 176.155 ;
    END
  END w_mask_in[1248]
  PIN w_mask_in[1249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.225 0.070 176.295 ;
    END
  END w_mask_in[1249]
  PIN w_mask_in[1250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.365 0.070 176.435 ;
    END
  END w_mask_in[1250]
  PIN w_mask_in[1251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.505 0.070 176.575 ;
    END
  END w_mask_in[1251]
  PIN w_mask_in[1252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.645 0.070 176.715 ;
    END
  END w_mask_in[1252]
  PIN w_mask_in[1253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.785 0.070 176.855 ;
    END
  END w_mask_in[1253]
  PIN w_mask_in[1254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.925 0.070 176.995 ;
    END
  END w_mask_in[1254]
  PIN w_mask_in[1255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.065 0.070 177.135 ;
    END
  END w_mask_in[1255]
  PIN w_mask_in[1256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.205 0.070 177.275 ;
    END
  END w_mask_in[1256]
  PIN w_mask_in[1257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.345 0.070 177.415 ;
    END
  END w_mask_in[1257]
  PIN w_mask_in[1258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.485 0.070 177.555 ;
    END
  END w_mask_in[1258]
  PIN w_mask_in[1259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.625 0.070 177.695 ;
    END
  END w_mask_in[1259]
  PIN w_mask_in[1260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END w_mask_in[1260]
  PIN w_mask_in[1261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.905 0.070 177.975 ;
    END
  END w_mask_in[1261]
  PIN w_mask_in[1262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.045 0.070 178.115 ;
    END
  END w_mask_in[1262]
  PIN w_mask_in[1263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.185 0.070 178.255 ;
    END
  END w_mask_in[1263]
  PIN w_mask_in[1264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.325 0.070 178.395 ;
    END
  END w_mask_in[1264]
  PIN w_mask_in[1265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.465 0.070 178.535 ;
    END
  END w_mask_in[1265]
  PIN w_mask_in[1266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.605 0.070 178.675 ;
    END
  END w_mask_in[1266]
  PIN w_mask_in[1267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.745 0.070 178.815 ;
    END
  END w_mask_in[1267]
  PIN w_mask_in[1268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.885 0.070 178.955 ;
    END
  END w_mask_in[1268]
  PIN w_mask_in[1269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.025 0.070 179.095 ;
    END
  END w_mask_in[1269]
  PIN w_mask_in[1270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.165 0.070 179.235 ;
    END
  END w_mask_in[1270]
  PIN w_mask_in[1271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.305 0.070 179.375 ;
    END
  END w_mask_in[1271]
  PIN w_mask_in[1272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.445 0.070 179.515 ;
    END
  END w_mask_in[1272]
  PIN w_mask_in[1273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.585 0.070 179.655 ;
    END
  END w_mask_in[1273]
  PIN w_mask_in[1274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END w_mask_in[1274]
  PIN w_mask_in[1275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.865 0.070 179.935 ;
    END
  END w_mask_in[1275]
  PIN w_mask_in[1276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.005 0.070 180.075 ;
    END
  END w_mask_in[1276]
  PIN w_mask_in[1277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.145 0.070 180.215 ;
    END
  END w_mask_in[1277]
  PIN w_mask_in[1278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.285 0.070 180.355 ;
    END
  END w_mask_in[1278]
  PIN w_mask_in[1279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.425 0.070 180.495 ;
    END
  END w_mask_in[1279]
  PIN w_mask_in[1280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.565 0.070 180.635 ;
    END
  END w_mask_in[1280]
  PIN w_mask_in[1281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.705 0.070 180.775 ;
    END
  END w_mask_in[1281]
  PIN w_mask_in[1282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.845 0.070 180.915 ;
    END
  END w_mask_in[1282]
  PIN w_mask_in[1283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.985 0.070 181.055 ;
    END
  END w_mask_in[1283]
  PIN w_mask_in[1284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.125 0.070 181.195 ;
    END
  END w_mask_in[1284]
  PIN w_mask_in[1285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.265 0.070 181.335 ;
    END
  END w_mask_in[1285]
  PIN w_mask_in[1286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.405 0.070 181.475 ;
    END
  END w_mask_in[1286]
  PIN w_mask_in[1287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.545 0.070 181.615 ;
    END
  END w_mask_in[1287]
  PIN w_mask_in[1288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.685 0.070 181.755 ;
    END
  END w_mask_in[1288]
  PIN w_mask_in[1289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.825 0.070 181.895 ;
    END
  END w_mask_in[1289]
  PIN w_mask_in[1290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.965 0.070 182.035 ;
    END
  END w_mask_in[1290]
  PIN w_mask_in[1291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.105 0.070 182.175 ;
    END
  END w_mask_in[1291]
  PIN w_mask_in[1292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.245 0.070 182.315 ;
    END
  END w_mask_in[1292]
  PIN w_mask_in[1293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.385 0.070 182.455 ;
    END
  END w_mask_in[1293]
  PIN w_mask_in[1294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.525 0.070 182.595 ;
    END
  END w_mask_in[1294]
  PIN w_mask_in[1295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.665 0.070 182.735 ;
    END
  END w_mask_in[1295]
  PIN w_mask_in[1296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.805 0.070 182.875 ;
    END
  END w_mask_in[1296]
  PIN w_mask_in[1297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.945 0.070 183.015 ;
    END
  END w_mask_in[1297]
  PIN w_mask_in[1298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.085 0.070 183.155 ;
    END
  END w_mask_in[1298]
  PIN w_mask_in[1299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.225 0.070 183.295 ;
    END
  END w_mask_in[1299]
  PIN w_mask_in[1300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.365 0.070 183.435 ;
    END
  END w_mask_in[1300]
  PIN w_mask_in[1301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.505 0.070 183.575 ;
    END
  END w_mask_in[1301]
  PIN w_mask_in[1302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.645 0.070 183.715 ;
    END
  END w_mask_in[1302]
  PIN w_mask_in[1303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.785 0.070 183.855 ;
    END
  END w_mask_in[1303]
  PIN w_mask_in[1304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.925 0.070 183.995 ;
    END
  END w_mask_in[1304]
  PIN w_mask_in[1305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.065 0.070 184.135 ;
    END
  END w_mask_in[1305]
  PIN w_mask_in[1306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.205 0.070 184.275 ;
    END
  END w_mask_in[1306]
  PIN w_mask_in[1307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.345 0.070 184.415 ;
    END
  END w_mask_in[1307]
  PIN w_mask_in[1308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.485 0.070 184.555 ;
    END
  END w_mask_in[1308]
  PIN w_mask_in[1309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.625 0.070 184.695 ;
    END
  END w_mask_in[1309]
  PIN w_mask_in[1310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.765 0.070 184.835 ;
    END
  END w_mask_in[1310]
  PIN w_mask_in[1311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.905 0.070 184.975 ;
    END
  END w_mask_in[1311]
  PIN w_mask_in[1312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.045 0.070 185.115 ;
    END
  END w_mask_in[1312]
  PIN w_mask_in[1313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.185 0.070 185.255 ;
    END
  END w_mask_in[1313]
  PIN w_mask_in[1314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.325 0.070 185.395 ;
    END
  END w_mask_in[1314]
  PIN w_mask_in[1315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.465 0.070 185.535 ;
    END
  END w_mask_in[1315]
  PIN w_mask_in[1316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.605 0.070 185.675 ;
    END
  END w_mask_in[1316]
  PIN w_mask_in[1317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.745 0.070 185.815 ;
    END
  END w_mask_in[1317]
  PIN w_mask_in[1318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.885 0.070 185.955 ;
    END
  END w_mask_in[1318]
  PIN w_mask_in[1319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.025 0.070 186.095 ;
    END
  END w_mask_in[1319]
  PIN w_mask_in[1320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.165 0.070 186.235 ;
    END
  END w_mask_in[1320]
  PIN w_mask_in[1321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.305 0.070 186.375 ;
    END
  END w_mask_in[1321]
  PIN w_mask_in[1322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.445 0.070 186.515 ;
    END
  END w_mask_in[1322]
  PIN w_mask_in[1323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.585 0.070 186.655 ;
    END
  END w_mask_in[1323]
  PIN w_mask_in[1324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.725 0.070 186.795 ;
    END
  END w_mask_in[1324]
  PIN w_mask_in[1325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.865 0.070 186.935 ;
    END
  END w_mask_in[1325]
  PIN w_mask_in[1326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.005 0.070 187.075 ;
    END
  END w_mask_in[1326]
  PIN w_mask_in[1327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.145 0.070 187.215 ;
    END
  END w_mask_in[1327]
  PIN w_mask_in[1328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.285 0.070 187.355 ;
    END
  END w_mask_in[1328]
  PIN w_mask_in[1329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.425 0.070 187.495 ;
    END
  END w_mask_in[1329]
  PIN w_mask_in[1330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.565 0.070 187.635 ;
    END
  END w_mask_in[1330]
  PIN w_mask_in[1331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.705 0.070 187.775 ;
    END
  END w_mask_in[1331]
  PIN w_mask_in[1332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.845 0.070 187.915 ;
    END
  END w_mask_in[1332]
  PIN w_mask_in[1333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.985 0.070 188.055 ;
    END
  END w_mask_in[1333]
  PIN w_mask_in[1334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END w_mask_in[1334]
  PIN w_mask_in[1335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.265 0.070 188.335 ;
    END
  END w_mask_in[1335]
  PIN w_mask_in[1336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.405 0.070 188.475 ;
    END
  END w_mask_in[1336]
  PIN w_mask_in[1337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.545 0.070 188.615 ;
    END
  END w_mask_in[1337]
  PIN w_mask_in[1338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.685 0.070 188.755 ;
    END
  END w_mask_in[1338]
  PIN w_mask_in[1339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.825 0.070 188.895 ;
    END
  END w_mask_in[1339]
  PIN w_mask_in[1340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.965 0.070 189.035 ;
    END
  END w_mask_in[1340]
  PIN w_mask_in[1341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.105 0.070 189.175 ;
    END
  END w_mask_in[1341]
  PIN w_mask_in[1342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.245 0.070 189.315 ;
    END
  END w_mask_in[1342]
  PIN w_mask_in[1343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.385 0.070 189.455 ;
    END
  END w_mask_in[1343]
  PIN w_mask_in[1344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.525 0.070 189.595 ;
    END
  END w_mask_in[1344]
  PIN w_mask_in[1345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.665 0.070 189.735 ;
    END
  END w_mask_in[1345]
  PIN w_mask_in[1346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.805 0.070 189.875 ;
    END
  END w_mask_in[1346]
  PIN w_mask_in[1347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.945 0.070 190.015 ;
    END
  END w_mask_in[1347]
  PIN w_mask_in[1348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.085 0.070 190.155 ;
    END
  END w_mask_in[1348]
  PIN w_mask_in[1349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.225 0.070 190.295 ;
    END
  END w_mask_in[1349]
  PIN w_mask_in[1350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.365 0.070 190.435 ;
    END
  END w_mask_in[1350]
  PIN w_mask_in[1351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.505 0.070 190.575 ;
    END
  END w_mask_in[1351]
  PIN w_mask_in[1352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.645 0.070 190.715 ;
    END
  END w_mask_in[1352]
  PIN w_mask_in[1353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.785 0.070 190.855 ;
    END
  END w_mask_in[1353]
  PIN w_mask_in[1354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.925 0.070 190.995 ;
    END
  END w_mask_in[1354]
  PIN w_mask_in[1355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.065 0.070 191.135 ;
    END
  END w_mask_in[1355]
  PIN w_mask_in[1356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.205 0.070 191.275 ;
    END
  END w_mask_in[1356]
  PIN w_mask_in[1357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.345 0.070 191.415 ;
    END
  END w_mask_in[1357]
  PIN w_mask_in[1358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.485 0.070 191.555 ;
    END
  END w_mask_in[1358]
  PIN w_mask_in[1359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.625 0.070 191.695 ;
    END
  END w_mask_in[1359]
  PIN w_mask_in[1360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.765 0.070 191.835 ;
    END
  END w_mask_in[1360]
  PIN w_mask_in[1361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.905 0.070 191.975 ;
    END
  END w_mask_in[1361]
  PIN w_mask_in[1362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.045 0.070 192.115 ;
    END
  END w_mask_in[1362]
  PIN w_mask_in[1363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.185 0.070 192.255 ;
    END
  END w_mask_in[1363]
  PIN w_mask_in[1364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.325 0.070 192.395 ;
    END
  END w_mask_in[1364]
  PIN w_mask_in[1365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.465 0.070 192.535 ;
    END
  END w_mask_in[1365]
  PIN w_mask_in[1366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.605 0.070 192.675 ;
    END
  END w_mask_in[1366]
  PIN w_mask_in[1367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.745 0.070 192.815 ;
    END
  END w_mask_in[1367]
  PIN w_mask_in[1368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.885 0.070 192.955 ;
    END
  END w_mask_in[1368]
  PIN w_mask_in[1369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.025 0.070 193.095 ;
    END
  END w_mask_in[1369]
  PIN w_mask_in[1370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.165 0.070 193.235 ;
    END
  END w_mask_in[1370]
  PIN w_mask_in[1371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.305 0.070 193.375 ;
    END
  END w_mask_in[1371]
  PIN w_mask_in[1372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.445 0.070 193.515 ;
    END
  END w_mask_in[1372]
  PIN w_mask_in[1373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.585 0.070 193.655 ;
    END
  END w_mask_in[1373]
  PIN w_mask_in[1374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.725 0.070 193.795 ;
    END
  END w_mask_in[1374]
  PIN w_mask_in[1375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.865 0.070 193.935 ;
    END
  END w_mask_in[1375]
  PIN w_mask_in[1376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.005 0.070 194.075 ;
    END
  END w_mask_in[1376]
  PIN w_mask_in[1377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.145 0.070 194.215 ;
    END
  END w_mask_in[1377]
  PIN w_mask_in[1378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.285 0.070 194.355 ;
    END
  END w_mask_in[1378]
  PIN w_mask_in[1379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.425 0.070 194.495 ;
    END
  END w_mask_in[1379]
  PIN w_mask_in[1380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.565 0.070 194.635 ;
    END
  END w_mask_in[1380]
  PIN w_mask_in[1381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.705 0.070 194.775 ;
    END
  END w_mask_in[1381]
  PIN w_mask_in[1382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.845 0.070 194.915 ;
    END
  END w_mask_in[1382]
  PIN w_mask_in[1383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.985 0.070 195.055 ;
    END
  END w_mask_in[1383]
  PIN w_mask_in[1384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.125 0.070 195.195 ;
    END
  END w_mask_in[1384]
  PIN w_mask_in[1385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.265 0.070 195.335 ;
    END
  END w_mask_in[1385]
  PIN w_mask_in[1386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.405 0.070 195.475 ;
    END
  END w_mask_in[1386]
  PIN w_mask_in[1387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.545 0.070 195.615 ;
    END
  END w_mask_in[1387]
  PIN w_mask_in[1388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.685 0.070 195.755 ;
    END
  END w_mask_in[1388]
  PIN w_mask_in[1389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.825 0.070 195.895 ;
    END
  END w_mask_in[1389]
  PIN w_mask_in[1390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.965 0.070 196.035 ;
    END
  END w_mask_in[1390]
  PIN w_mask_in[1391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.105 0.070 196.175 ;
    END
  END w_mask_in[1391]
  PIN w_mask_in[1392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.245 0.070 196.315 ;
    END
  END w_mask_in[1392]
  PIN w_mask_in[1393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.385 0.070 196.455 ;
    END
  END w_mask_in[1393]
  PIN w_mask_in[1394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.525 0.070 196.595 ;
    END
  END w_mask_in[1394]
  PIN w_mask_in[1395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.665 0.070 196.735 ;
    END
  END w_mask_in[1395]
  PIN w_mask_in[1396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.805 0.070 196.875 ;
    END
  END w_mask_in[1396]
  PIN w_mask_in[1397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.945 0.070 197.015 ;
    END
  END w_mask_in[1397]
  PIN w_mask_in[1398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.085 0.070 197.155 ;
    END
  END w_mask_in[1398]
  PIN w_mask_in[1399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.225 0.070 197.295 ;
    END
  END w_mask_in[1399]
  PIN w_mask_in[1400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END w_mask_in[1400]
  PIN w_mask_in[1401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.505 0.070 197.575 ;
    END
  END w_mask_in[1401]
  PIN w_mask_in[1402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.645 0.070 197.715 ;
    END
  END w_mask_in[1402]
  PIN w_mask_in[1403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.785 0.070 197.855 ;
    END
  END w_mask_in[1403]
  PIN w_mask_in[1404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.925 0.070 197.995 ;
    END
  END w_mask_in[1404]
  PIN w_mask_in[1405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.065 0.070 198.135 ;
    END
  END w_mask_in[1405]
  PIN w_mask_in[1406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.205 0.070 198.275 ;
    END
  END w_mask_in[1406]
  PIN w_mask_in[1407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.345 0.070 198.415 ;
    END
  END w_mask_in[1407]
  PIN w_mask_in[1408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.485 0.070 198.555 ;
    END
  END w_mask_in[1408]
  PIN w_mask_in[1409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.625 0.070 198.695 ;
    END
  END w_mask_in[1409]
  PIN w_mask_in[1410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.765 0.070 198.835 ;
    END
  END w_mask_in[1410]
  PIN w_mask_in[1411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.905 0.070 198.975 ;
    END
  END w_mask_in[1411]
  PIN w_mask_in[1412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.045 0.070 199.115 ;
    END
  END w_mask_in[1412]
  PIN w_mask_in[1413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.185 0.070 199.255 ;
    END
  END w_mask_in[1413]
  PIN w_mask_in[1414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.325 0.070 199.395 ;
    END
  END w_mask_in[1414]
  PIN w_mask_in[1415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.465 0.070 199.535 ;
    END
  END w_mask_in[1415]
  PIN w_mask_in[1416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.605 0.070 199.675 ;
    END
  END w_mask_in[1416]
  PIN w_mask_in[1417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.745 0.070 199.815 ;
    END
  END w_mask_in[1417]
  PIN w_mask_in[1418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.885 0.070 199.955 ;
    END
  END w_mask_in[1418]
  PIN w_mask_in[1419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.025 0.070 200.095 ;
    END
  END w_mask_in[1419]
  PIN w_mask_in[1420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.165 0.070 200.235 ;
    END
  END w_mask_in[1420]
  PIN w_mask_in[1421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.305 0.070 200.375 ;
    END
  END w_mask_in[1421]
  PIN w_mask_in[1422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.445 0.070 200.515 ;
    END
  END w_mask_in[1422]
  PIN w_mask_in[1423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.585 0.070 200.655 ;
    END
  END w_mask_in[1423]
  PIN w_mask_in[1424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.725 0.070 200.795 ;
    END
  END w_mask_in[1424]
  PIN w_mask_in[1425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.865 0.070 200.935 ;
    END
  END w_mask_in[1425]
  PIN w_mask_in[1426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.005 0.070 201.075 ;
    END
  END w_mask_in[1426]
  PIN w_mask_in[1427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.145 0.070 201.215 ;
    END
  END w_mask_in[1427]
  PIN w_mask_in[1428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.285 0.070 201.355 ;
    END
  END w_mask_in[1428]
  PIN w_mask_in[1429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.425 0.070 201.495 ;
    END
  END w_mask_in[1429]
  PIN w_mask_in[1430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.565 0.070 201.635 ;
    END
  END w_mask_in[1430]
  PIN w_mask_in[1431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.705 0.070 201.775 ;
    END
  END w_mask_in[1431]
  PIN w_mask_in[1432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.845 0.070 201.915 ;
    END
  END w_mask_in[1432]
  PIN w_mask_in[1433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.985 0.070 202.055 ;
    END
  END w_mask_in[1433]
  PIN w_mask_in[1434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.125 0.070 202.195 ;
    END
  END w_mask_in[1434]
  PIN w_mask_in[1435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.265 0.070 202.335 ;
    END
  END w_mask_in[1435]
  PIN w_mask_in[1436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.405 0.070 202.475 ;
    END
  END w_mask_in[1436]
  PIN w_mask_in[1437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.545 0.070 202.615 ;
    END
  END w_mask_in[1437]
  PIN w_mask_in[1438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.685 0.070 202.755 ;
    END
  END w_mask_in[1438]
  PIN w_mask_in[1439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.825 0.070 202.895 ;
    END
  END w_mask_in[1439]
  PIN w_mask_in[1440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.965 0.070 203.035 ;
    END
  END w_mask_in[1440]
  PIN w_mask_in[1441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.105 0.070 203.175 ;
    END
  END w_mask_in[1441]
  PIN w_mask_in[1442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.245 0.070 203.315 ;
    END
  END w_mask_in[1442]
  PIN w_mask_in[1443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.385 0.070 203.455 ;
    END
  END w_mask_in[1443]
  PIN w_mask_in[1444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.525 0.070 203.595 ;
    END
  END w_mask_in[1444]
  PIN w_mask_in[1445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.665 0.070 203.735 ;
    END
  END w_mask_in[1445]
  PIN w_mask_in[1446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.805 0.070 203.875 ;
    END
  END w_mask_in[1446]
  PIN w_mask_in[1447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.945 0.070 204.015 ;
    END
  END w_mask_in[1447]
  PIN w_mask_in[1448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.085 0.070 204.155 ;
    END
  END w_mask_in[1448]
  PIN w_mask_in[1449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.225 0.070 204.295 ;
    END
  END w_mask_in[1449]
  PIN w_mask_in[1450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.365 0.070 204.435 ;
    END
  END w_mask_in[1450]
  PIN w_mask_in[1451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.505 0.070 204.575 ;
    END
  END w_mask_in[1451]
  PIN w_mask_in[1452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.645 0.070 204.715 ;
    END
  END w_mask_in[1452]
  PIN w_mask_in[1453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.785 0.070 204.855 ;
    END
  END w_mask_in[1453]
  PIN w_mask_in[1454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.925 0.070 204.995 ;
    END
  END w_mask_in[1454]
  PIN w_mask_in[1455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.065 0.070 205.135 ;
    END
  END w_mask_in[1455]
  PIN w_mask_in[1456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.205 0.070 205.275 ;
    END
  END w_mask_in[1456]
  PIN w_mask_in[1457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.345 0.070 205.415 ;
    END
  END w_mask_in[1457]
  PIN w_mask_in[1458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.485 0.070 205.555 ;
    END
  END w_mask_in[1458]
  PIN w_mask_in[1459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.625 0.070 205.695 ;
    END
  END w_mask_in[1459]
  PIN w_mask_in[1460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.765 0.070 205.835 ;
    END
  END w_mask_in[1460]
  PIN w_mask_in[1461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.905 0.070 205.975 ;
    END
  END w_mask_in[1461]
  PIN w_mask_in[1462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.045 0.070 206.115 ;
    END
  END w_mask_in[1462]
  PIN w_mask_in[1463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.185 0.070 206.255 ;
    END
  END w_mask_in[1463]
  PIN w_mask_in[1464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.325 0.070 206.395 ;
    END
  END w_mask_in[1464]
  PIN w_mask_in[1465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.465 0.070 206.535 ;
    END
  END w_mask_in[1465]
  PIN w_mask_in[1466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.605 0.070 206.675 ;
    END
  END w_mask_in[1466]
  PIN w_mask_in[1467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.745 0.070 206.815 ;
    END
  END w_mask_in[1467]
  PIN w_mask_in[1468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.885 0.070 206.955 ;
    END
  END w_mask_in[1468]
  PIN w_mask_in[1469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.025 0.070 207.095 ;
    END
  END w_mask_in[1469]
  PIN w_mask_in[1470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.165 0.070 207.235 ;
    END
  END w_mask_in[1470]
  PIN w_mask_in[1471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.305 0.070 207.375 ;
    END
  END w_mask_in[1471]
  PIN w_mask_in[1472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.445 0.070 207.515 ;
    END
  END w_mask_in[1472]
  PIN w_mask_in[1473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.585 0.070 207.655 ;
    END
  END w_mask_in[1473]
  PIN w_mask_in[1474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.725 0.070 207.795 ;
    END
  END w_mask_in[1474]
  PIN w_mask_in[1475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.865 0.070 207.935 ;
    END
  END w_mask_in[1475]
  PIN w_mask_in[1476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.005 0.070 208.075 ;
    END
  END w_mask_in[1476]
  PIN w_mask_in[1477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.145 0.070 208.215 ;
    END
  END w_mask_in[1477]
  PIN w_mask_in[1478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.285 0.070 208.355 ;
    END
  END w_mask_in[1478]
  PIN w_mask_in[1479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.425 0.070 208.495 ;
    END
  END w_mask_in[1479]
  PIN w_mask_in[1480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.565 0.070 208.635 ;
    END
  END w_mask_in[1480]
  PIN w_mask_in[1481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.705 0.070 208.775 ;
    END
  END w_mask_in[1481]
  PIN w_mask_in[1482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.845 0.070 208.915 ;
    END
  END w_mask_in[1482]
  PIN w_mask_in[1483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.985 0.070 209.055 ;
    END
  END w_mask_in[1483]
  PIN w_mask_in[1484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.125 0.070 209.195 ;
    END
  END w_mask_in[1484]
  PIN w_mask_in[1485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.265 0.070 209.335 ;
    END
  END w_mask_in[1485]
  PIN w_mask_in[1486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.405 0.070 209.475 ;
    END
  END w_mask_in[1486]
  PIN w_mask_in[1487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.545 0.070 209.615 ;
    END
  END w_mask_in[1487]
  PIN w_mask_in[1488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.685 0.070 209.755 ;
    END
  END w_mask_in[1488]
  PIN w_mask_in[1489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.825 0.070 209.895 ;
    END
  END w_mask_in[1489]
  PIN w_mask_in[1490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.965 0.070 210.035 ;
    END
  END w_mask_in[1490]
  PIN w_mask_in[1491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.105 0.070 210.175 ;
    END
  END w_mask_in[1491]
  PIN w_mask_in[1492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.245 0.070 210.315 ;
    END
  END w_mask_in[1492]
  PIN w_mask_in[1493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.385 0.070 210.455 ;
    END
  END w_mask_in[1493]
  PIN w_mask_in[1494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END w_mask_in[1494]
  PIN w_mask_in[1495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.665 0.070 210.735 ;
    END
  END w_mask_in[1495]
  PIN w_mask_in[1496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.805 0.070 210.875 ;
    END
  END w_mask_in[1496]
  PIN w_mask_in[1497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.945 0.070 211.015 ;
    END
  END w_mask_in[1497]
  PIN w_mask_in[1498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.085 0.070 211.155 ;
    END
  END w_mask_in[1498]
  PIN w_mask_in[1499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.225 0.070 211.295 ;
    END
  END w_mask_in[1499]
  PIN w_mask_in[1500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.365 0.070 211.435 ;
    END
  END w_mask_in[1500]
  PIN w_mask_in[1501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.505 0.070 211.575 ;
    END
  END w_mask_in[1501]
  PIN w_mask_in[1502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.645 0.070 211.715 ;
    END
  END w_mask_in[1502]
  PIN w_mask_in[1503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.785 0.070 211.855 ;
    END
  END w_mask_in[1503]
  PIN w_mask_in[1504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 211.925 0.070 211.995 ;
    END
  END w_mask_in[1504]
  PIN w_mask_in[1505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.065 0.070 212.135 ;
    END
  END w_mask_in[1505]
  PIN w_mask_in[1506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.205 0.070 212.275 ;
    END
  END w_mask_in[1506]
  PIN w_mask_in[1507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.345 0.070 212.415 ;
    END
  END w_mask_in[1507]
  PIN w_mask_in[1508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.485 0.070 212.555 ;
    END
  END w_mask_in[1508]
  PIN w_mask_in[1509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.625 0.070 212.695 ;
    END
  END w_mask_in[1509]
  PIN w_mask_in[1510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.765 0.070 212.835 ;
    END
  END w_mask_in[1510]
  PIN w_mask_in[1511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.905 0.070 212.975 ;
    END
  END w_mask_in[1511]
  PIN w_mask_in[1512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.045 0.070 213.115 ;
    END
  END w_mask_in[1512]
  PIN w_mask_in[1513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.185 0.070 213.255 ;
    END
  END w_mask_in[1513]
  PIN w_mask_in[1514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.325 0.070 213.395 ;
    END
  END w_mask_in[1514]
  PIN w_mask_in[1515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.465 0.070 213.535 ;
    END
  END w_mask_in[1515]
  PIN w_mask_in[1516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.605 0.070 213.675 ;
    END
  END w_mask_in[1516]
  PIN w_mask_in[1517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.745 0.070 213.815 ;
    END
  END w_mask_in[1517]
  PIN w_mask_in[1518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.885 0.070 213.955 ;
    END
  END w_mask_in[1518]
  PIN w_mask_in[1519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.025 0.070 214.095 ;
    END
  END w_mask_in[1519]
  PIN w_mask_in[1520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.165 0.070 214.235 ;
    END
  END w_mask_in[1520]
  PIN w_mask_in[1521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.305 0.070 214.375 ;
    END
  END w_mask_in[1521]
  PIN w_mask_in[1522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.445 0.070 214.515 ;
    END
  END w_mask_in[1522]
  PIN w_mask_in[1523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.585 0.070 214.655 ;
    END
  END w_mask_in[1523]
  PIN w_mask_in[1524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.725 0.070 214.795 ;
    END
  END w_mask_in[1524]
  PIN w_mask_in[1525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 214.865 0.070 214.935 ;
    END
  END w_mask_in[1525]
  PIN w_mask_in[1526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END w_mask_in[1526]
  PIN w_mask_in[1527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.145 0.070 215.215 ;
    END
  END w_mask_in[1527]
  PIN w_mask_in[1528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.285 0.070 215.355 ;
    END
  END w_mask_in[1528]
  PIN w_mask_in[1529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.425 0.070 215.495 ;
    END
  END w_mask_in[1529]
  PIN w_mask_in[1530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.565 0.070 215.635 ;
    END
  END w_mask_in[1530]
  PIN w_mask_in[1531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.705 0.070 215.775 ;
    END
  END w_mask_in[1531]
  PIN w_mask_in[1532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.845 0.070 215.915 ;
    END
  END w_mask_in[1532]
  PIN w_mask_in[1533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.985 0.070 216.055 ;
    END
  END w_mask_in[1533]
  PIN w_mask_in[1534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.125 0.070 216.195 ;
    END
  END w_mask_in[1534]
  PIN w_mask_in[1535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.265 0.070 216.335 ;
    END
  END w_mask_in[1535]
  PIN w_mask_in[1536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.405 0.070 216.475 ;
    END
  END w_mask_in[1536]
  PIN w_mask_in[1537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.545 0.070 216.615 ;
    END
  END w_mask_in[1537]
  PIN w_mask_in[1538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.685 0.070 216.755 ;
    END
  END w_mask_in[1538]
  PIN w_mask_in[1539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.825 0.070 216.895 ;
    END
  END w_mask_in[1539]
  PIN w_mask_in[1540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.965 0.070 217.035 ;
    END
  END w_mask_in[1540]
  PIN w_mask_in[1541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.105 0.070 217.175 ;
    END
  END w_mask_in[1541]
  PIN w_mask_in[1542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.245 0.070 217.315 ;
    END
  END w_mask_in[1542]
  PIN w_mask_in[1543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.385 0.070 217.455 ;
    END
  END w_mask_in[1543]
  PIN w_mask_in[1544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.525 0.070 217.595 ;
    END
  END w_mask_in[1544]
  PIN w_mask_in[1545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.665 0.070 217.735 ;
    END
  END w_mask_in[1545]
  PIN w_mask_in[1546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.805 0.070 217.875 ;
    END
  END w_mask_in[1546]
  PIN w_mask_in[1547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.945 0.070 218.015 ;
    END
  END w_mask_in[1547]
  PIN w_mask_in[1548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.085 0.070 218.155 ;
    END
  END w_mask_in[1548]
  PIN w_mask_in[1549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.225 0.070 218.295 ;
    END
  END w_mask_in[1549]
  PIN w_mask_in[1550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.365 0.070 218.435 ;
    END
  END w_mask_in[1550]
  PIN w_mask_in[1551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.505 0.070 218.575 ;
    END
  END w_mask_in[1551]
  PIN w_mask_in[1552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.645 0.070 218.715 ;
    END
  END w_mask_in[1552]
  PIN w_mask_in[1553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.785 0.070 218.855 ;
    END
  END w_mask_in[1553]
  PIN w_mask_in[1554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.925 0.070 218.995 ;
    END
  END w_mask_in[1554]
  PIN w_mask_in[1555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.065 0.070 219.135 ;
    END
  END w_mask_in[1555]
  PIN w_mask_in[1556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.205 0.070 219.275 ;
    END
  END w_mask_in[1556]
  PIN w_mask_in[1557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.345 0.070 219.415 ;
    END
  END w_mask_in[1557]
  PIN w_mask_in[1558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.485 0.070 219.555 ;
    END
  END w_mask_in[1558]
  PIN w_mask_in[1559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.625 0.070 219.695 ;
    END
  END w_mask_in[1559]
  PIN w_mask_in[1560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.765 0.070 219.835 ;
    END
  END w_mask_in[1560]
  PIN w_mask_in[1561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 219.905 0.070 219.975 ;
    END
  END w_mask_in[1561]
  PIN w_mask_in[1562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.045 0.070 220.115 ;
    END
  END w_mask_in[1562]
  PIN w_mask_in[1563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.185 0.070 220.255 ;
    END
  END w_mask_in[1563]
  PIN w_mask_in[1564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.325 0.070 220.395 ;
    END
  END w_mask_in[1564]
  PIN w_mask_in[1565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.465 0.070 220.535 ;
    END
  END w_mask_in[1565]
  PIN w_mask_in[1566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.605 0.070 220.675 ;
    END
  END w_mask_in[1566]
  PIN w_mask_in[1567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.745 0.070 220.815 ;
    END
  END w_mask_in[1567]
  PIN w_mask_in[1568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.885 0.070 220.955 ;
    END
  END w_mask_in[1568]
  PIN w_mask_in[1569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.025 0.070 221.095 ;
    END
  END w_mask_in[1569]
  PIN w_mask_in[1570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.165 0.070 221.235 ;
    END
  END w_mask_in[1570]
  PIN w_mask_in[1571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.305 0.070 221.375 ;
    END
  END w_mask_in[1571]
  PIN w_mask_in[1572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.445 0.070 221.515 ;
    END
  END w_mask_in[1572]
  PIN w_mask_in[1573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.585 0.070 221.655 ;
    END
  END w_mask_in[1573]
  PIN w_mask_in[1574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.725 0.070 221.795 ;
    END
  END w_mask_in[1574]
  PIN w_mask_in[1575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.865 0.070 221.935 ;
    END
  END w_mask_in[1575]
  PIN w_mask_in[1576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.005 0.070 222.075 ;
    END
  END w_mask_in[1576]
  PIN w_mask_in[1577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.145 0.070 222.215 ;
    END
  END w_mask_in[1577]
  PIN w_mask_in[1578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.285 0.070 222.355 ;
    END
  END w_mask_in[1578]
  PIN w_mask_in[1579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.425 0.070 222.495 ;
    END
  END w_mask_in[1579]
  PIN w_mask_in[1580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.565 0.070 222.635 ;
    END
  END w_mask_in[1580]
  PIN w_mask_in[1581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.705 0.070 222.775 ;
    END
  END w_mask_in[1581]
  PIN w_mask_in[1582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.845 0.070 222.915 ;
    END
  END w_mask_in[1582]
  PIN w_mask_in[1583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 222.985 0.070 223.055 ;
    END
  END w_mask_in[1583]
  PIN w_mask_in[1584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.125 0.070 223.195 ;
    END
  END w_mask_in[1584]
  PIN w_mask_in[1585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.265 0.070 223.335 ;
    END
  END w_mask_in[1585]
  PIN w_mask_in[1586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.405 0.070 223.475 ;
    END
  END w_mask_in[1586]
  PIN w_mask_in[1587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.545 0.070 223.615 ;
    END
  END w_mask_in[1587]
  PIN w_mask_in[1588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.685 0.070 223.755 ;
    END
  END w_mask_in[1588]
  PIN w_mask_in[1589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.825 0.070 223.895 ;
    END
  END w_mask_in[1589]
  PIN w_mask_in[1590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.965 0.070 224.035 ;
    END
  END w_mask_in[1590]
  PIN w_mask_in[1591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.105 0.070 224.175 ;
    END
  END w_mask_in[1591]
  PIN w_mask_in[1592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.245 0.070 224.315 ;
    END
  END w_mask_in[1592]
  PIN w_mask_in[1593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.385 0.070 224.455 ;
    END
  END w_mask_in[1593]
  PIN w_mask_in[1594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.525 0.070 224.595 ;
    END
  END w_mask_in[1594]
  PIN w_mask_in[1595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.665 0.070 224.735 ;
    END
  END w_mask_in[1595]
  PIN w_mask_in[1596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.805 0.070 224.875 ;
    END
  END w_mask_in[1596]
  PIN w_mask_in[1597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.945 0.070 225.015 ;
    END
  END w_mask_in[1597]
  PIN w_mask_in[1598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.085 0.070 225.155 ;
    END
  END w_mask_in[1598]
  PIN w_mask_in[1599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.225 0.070 225.295 ;
    END
  END w_mask_in[1599]
  PIN w_mask_in[1600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.365 0.070 225.435 ;
    END
  END w_mask_in[1600]
  PIN w_mask_in[1601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.505 0.070 225.575 ;
    END
  END w_mask_in[1601]
  PIN w_mask_in[1602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.645 0.070 225.715 ;
    END
  END w_mask_in[1602]
  PIN w_mask_in[1603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.785 0.070 225.855 ;
    END
  END w_mask_in[1603]
  PIN w_mask_in[1604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 225.925 0.070 225.995 ;
    END
  END w_mask_in[1604]
  PIN w_mask_in[1605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.065 0.070 226.135 ;
    END
  END w_mask_in[1605]
  PIN w_mask_in[1606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.205 0.070 226.275 ;
    END
  END w_mask_in[1606]
  PIN w_mask_in[1607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.345 0.070 226.415 ;
    END
  END w_mask_in[1607]
  PIN w_mask_in[1608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.485 0.070 226.555 ;
    END
  END w_mask_in[1608]
  PIN w_mask_in[1609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.625 0.070 226.695 ;
    END
  END w_mask_in[1609]
  PIN w_mask_in[1610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END w_mask_in[1610]
  PIN w_mask_in[1611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.905 0.070 226.975 ;
    END
  END w_mask_in[1611]
  PIN w_mask_in[1612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.045 0.070 227.115 ;
    END
  END w_mask_in[1612]
  PIN w_mask_in[1613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.185 0.070 227.255 ;
    END
  END w_mask_in[1613]
  PIN w_mask_in[1614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.325 0.070 227.395 ;
    END
  END w_mask_in[1614]
  PIN w_mask_in[1615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.465 0.070 227.535 ;
    END
  END w_mask_in[1615]
  PIN w_mask_in[1616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.605 0.070 227.675 ;
    END
  END w_mask_in[1616]
  PIN w_mask_in[1617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.745 0.070 227.815 ;
    END
  END w_mask_in[1617]
  PIN w_mask_in[1618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.885 0.070 227.955 ;
    END
  END w_mask_in[1618]
  PIN w_mask_in[1619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.025 0.070 228.095 ;
    END
  END w_mask_in[1619]
  PIN w_mask_in[1620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.165 0.070 228.235 ;
    END
  END w_mask_in[1620]
  PIN w_mask_in[1621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.305 0.070 228.375 ;
    END
  END w_mask_in[1621]
  PIN w_mask_in[1622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.445 0.070 228.515 ;
    END
  END w_mask_in[1622]
  PIN w_mask_in[1623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.585 0.070 228.655 ;
    END
  END w_mask_in[1623]
  PIN w_mask_in[1624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.725 0.070 228.795 ;
    END
  END w_mask_in[1624]
  PIN w_mask_in[1625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 228.865 0.070 228.935 ;
    END
  END w_mask_in[1625]
  PIN w_mask_in[1626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.005 0.070 229.075 ;
    END
  END w_mask_in[1626]
  PIN w_mask_in[1627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.145 0.070 229.215 ;
    END
  END w_mask_in[1627]
  PIN w_mask_in[1628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.285 0.070 229.355 ;
    END
  END w_mask_in[1628]
  PIN w_mask_in[1629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.425 0.070 229.495 ;
    END
  END w_mask_in[1629]
  PIN w_mask_in[1630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.565 0.070 229.635 ;
    END
  END w_mask_in[1630]
  PIN w_mask_in[1631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.705 0.070 229.775 ;
    END
  END w_mask_in[1631]
  PIN w_mask_in[1632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.845 0.070 229.915 ;
    END
  END w_mask_in[1632]
  PIN w_mask_in[1633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.985 0.070 230.055 ;
    END
  END w_mask_in[1633]
  PIN w_mask_in[1634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.125 0.070 230.195 ;
    END
  END w_mask_in[1634]
  PIN w_mask_in[1635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.265 0.070 230.335 ;
    END
  END w_mask_in[1635]
  PIN w_mask_in[1636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.405 0.070 230.475 ;
    END
  END w_mask_in[1636]
  PIN w_mask_in[1637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.545 0.070 230.615 ;
    END
  END w_mask_in[1637]
  PIN w_mask_in[1638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.685 0.070 230.755 ;
    END
  END w_mask_in[1638]
  PIN w_mask_in[1639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.825 0.070 230.895 ;
    END
  END w_mask_in[1639]
  PIN w_mask_in[1640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.965 0.070 231.035 ;
    END
  END w_mask_in[1640]
  PIN w_mask_in[1641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.105 0.070 231.175 ;
    END
  END w_mask_in[1641]
  PIN w_mask_in[1642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.245 0.070 231.315 ;
    END
  END w_mask_in[1642]
  PIN w_mask_in[1643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.385 0.070 231.455 ;
    END
  END w_mask_in[1643]
  PIN w_mask_in[1644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.525 0.070 231.595 ;
    END
  END w_mask_in[1644]
  PIN w_mask_in[1645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.665 0.070 231.735 ;
    END
  END w_mask_in[1645]
  PIN w_mask_in[1646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.805 0.070 231.875 ;
    END
  END w_mask_in[1646]
  PIN w_mask_in[1647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.945 0.070 232.015 ;
    END
  END w_mask_in[1647]
  PIN w_mask_in[1648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.085 0.070 232.155 ;
    END
  END w_mask_in[1648]
  PIN w_mask_in[1649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.225 0.070 232.295 ;
    END
  END w_mask_in[1649]
  PIN w_mask_in[1650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.365 0.070 232.435 ;
    END
  END w_mask_in[1650]
  PIN w_mask_in[1651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.505 0.070 232.575 ;
    END
  END w_mask_in[1651]
  PIN w_mask_in[1652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.645 0.070 232.715 ;
    END
  END w_mask_in[1652]
  PIN w_mask_in[1653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.785 0.070 232.855 ;
    END
  END w_mask_in[1653]
  PIN w_mask_in[1654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.925 0.070 232.995 ;
    END
  END w_mask_in[1654]
  PIN w_mask_in[1655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.065 0.070 233.135 ;
    END
  END w_mask_in[1655]
  PIN w_mask_in[1656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.205 0.070 233.275 ;
    END
  END w_mask_in[1656]
  PIN w_mask_in[1657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.345 0.070 233.415 ;
    END
  END w_mask_in[1657]
  PIN w_mask_in[1658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.485 0.070 233.555 ;
    END
  END w_mask_in[1658]
  PIN w_mask_in[1659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.625 0.070 233.695 ;
    END
  END w_mask_in[1659]
  PIN w_mask_in[1660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.765 0.070 233.835 ;
    END
  END w_mask_in[1660]
  PIN w_mask_in[1661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.905 0.070 233.975 ;
    END
  END w_mask_in[1661]
  PIN w_mask_in[1662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.045 0.070 234.115 ;
    END
  END w_mask_in[1662]
  PIN w_mask_in[1663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.185 0.070 234.255 ;
    END
  END w_mask_in[1663]
  PIN w_mask_in[1664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.325 0.070 234.395 ;
    END
  END w_mask_in[1664]
  PIN w_mask_in[1665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.465 0.070 234.535 ;
    END
  END w_mask_in[1665]
  PIN w_mask_in[1666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.605 0.070 234.675 ;
    END
  END w_mask_in[1666]
  PIN w_mask_in[1667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.745 0.070 234.815 ;
    END
  END w_mask_in[1667]
  PIN w_mask_in[1668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.885 0.070 234.955 ;
    END
  END w_mask_in[1668]
  PIN w_mask_in[1669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.025 0.070 235.095 ;
    END
  END w_mask_in[1669]
  PIN w_mask_in[1670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.165 0.070 235.235 ;
    END
  END w_mask_in[1670]
  PIN w_mask_in[1671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.305 0.070 235.375 ;
    END
  END w_mask_in[1671]
  PIN w_mask_in[1672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.445 0.070 235.515 ;
    END
  END w_mask_in[1672]
  PIN w_mask_in[1673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.585 0.070 235.655 ;
    END
  END w_mask_in[1673]
  PIN w_mask_in[1674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.725 0.070 235.795 ;
    END
  END w_mask_in[1674]
  PIN w_mask_in[1675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.865 0.070 235.935 ;
    END
  END w_mask_in[1675]
  PIN w_mask_in[1676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.005 0.070 236.075 ;
    END
  END w_mask_in[1676]
  PIN w_mask_in[1677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.145 0.070 236.215 ;
    END
  END w_mask_in[1677]
  PIN w_mask_in[1678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.285 0.070 236.355 ;
    END
  END w_mask_in[1678]
  PIN w_mask_in[1679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.425 0.070 236.495 ;
    END
  END w_mask_in[1679]
  PIN w_mask_in[1680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.565 0.070 236.635 ;
    END
  END w_mask_in[1680]
  PIN w_mask_in[1681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.705 0.070 236.775 ;
    END
  END w_mask_in[1681]
  PIN w_mask_in[1682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.845 0.070 236.915 ;
    END
  END w_mask_in[1682]
  PIN w_mask_in[1683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.985 0.070 237.055 ;
    END
  END w_mask_in[1683]
  PIN w_mask_in[1684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.125 0.070 237.195 ;
    END
  END w_mask_in[1684]
  PIN w_mask_in[1685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.265 0.070 237.335 ;
    END
  END w_mask_in[1685]
  PIN w_mask_in[1686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.405 0.070 237.475 ;
    END
  END w_mask_in[1686]
  PIN w_mask_in[1687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.545 0.070 237.615 ;
    END
  END w_mask_in[1687]
  PIN w_mask_in[1688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.685 0.070 237.755 ;
    END
  END w_mask_in[1688]
  PIN w_mask_in[1689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.825 0.070 237.895 ;
    END
  END w_mask_in[1689]
  PIN w_mask_in[1690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 237.965 0.070 238.035 ;
    END
  END w_mask_in[1690]
  PIN w_mask_in[1691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.105 0.070 238.175 ;
    END
  END w_mask_in[1691]
  PIN w_mask_in[1692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.245 0.070 238.315 ;
    END
  END w_mask_in[1692]
  PIN w_mask_in[1693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.385 0.070 238.455 ;
    END
  END w_mask_in[1693]
  PIN w_mask_in[1694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.525 0.070 238.595 ;
    END
  END w_mask_in[1694]
  PIN w_mask_in[1695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.665 0.070 238.735 ;
    END
  END w_mask_in[1695]
  PIN w_mask_in[1696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.805 0.070 238.875 ;
    END
  END w_mask_in[1696]
  PIN w_mask_in[1697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.945 0.070 239.015 ;
    END
  END w_mask_in[1697]
  PIN w_mask_in[1698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.085 0.070 239.155 ;
    END
  END w_mask_in[1698]
  PIN w_mask_in[1699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.225 0.070 239.295 ;
    END
  END w_mask_in[1699]
  PIN w_mask_in[1700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.365 0.070 239.435 ;
    END
  END w_mask_in[1700]
  PIN w_mask_in[1701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.505 0.070 239.575 ;
    END
  END w_mask_in[1701]
  PIN w_mask_in[1702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.645 0.070 239.715 ;
    END
  END w_mask_in[1702]
  PIN w_mask_in[1703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.785 0.070 239.855 ;
    END
  END w_mask_in[1703]
  PIN w_mask_in[1704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.925 0.070 239.995 ;
    END
  END w_mask_in[1704]
  PIN w_mask_in[1705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.065 0.070 240.135 ;
    END
  END w_mask_in[1705]
  PIN w_mask_in[1706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.205 0.070 240.275 ;
    END
  END w_mask_in[1706]
  PIN w_mask_in[1707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.345 0.070 240.415 ;
    END
  END w_mask_in[1707]
  PIN w_mask_in[1708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.485 0.070 240.555 ;
    END
  END w_mask_in[1708]
  PIN w_mask_in[1709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.625 0.070 240.695 ;
    END
  END w_mask_in[1709]
  PIN w_mask_in[1710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.765 0.070 240.835 ;
    END
  END w_mask_in[1710]
  PIN w_mask_in[1711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 240.905 0.070 240.975 ;
    END
  END w_mask_in[1711]
  PIN w_mask_in[1712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.045 0.070 241.115 ;
    END
  END w_mask_in[1712]
  PIN w_mask_in[1713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.185 0.070 241.255 ;
    END
  END w_mask_in[1713]
  PIN w_mask_in[1714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.325 0.070 241.395 ;
    END
  END w_mask_in[1714]
  PIN w_mask_in[1715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.465 0.070 241.535 ;
    END
  END w_mask_in[1715]
  PIN w_mask_in[1716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.605 0.070 241.675 ;
    END
  END w_mask_in[1716]
  PIN w_mask_in[1717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.745 0.070 241.815 ;
    END
  END w_mask_in[1717]
  PIN w_mask_in[1718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.885 0.070 241.955 ;
    END
  END w_mask_in[1718]
  PIN w_mask_in[1719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.025 0.070 242.095 ;
    END
  END w_mask_in[1719]
  PIN w_mask_in[1720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.165 0.070 242.235 ;
    END
  END w_mask_in[1720]
  PIN w_mask_in[1721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.305 0.070 242.375 ;
    END
  END w_mask_in[1721]
  PIN w_mask_in[1722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.445 0.070 242.515 ;
    END
  END w_mask_in[1722]
  PIN w_mask_in[1723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.585 0.070 242.655 ;
    END
  END w_mask_in[1723]
  PIN w_mask_in[1724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.725 0.070 242.795 ;
    END
  END w_mask_in[1724]
  PIN w_mask_in[1725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 242.865 0.070 242.935 ;
    END
  END w_mask_in[1725]
  PIN w_mask_in[1726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.005 0.070 243.075 ;
    END
  END w_mask_in[1726]
  PIN w_mask_in[1727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.145 0.070 243.215 ;
    END
  END w_mask_in[1727]
  PIN w_mask_in[1728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.285 0.070 243.355 ;
    END
  END w_mask_in[1728]
  PIN w_mask_in[1729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.425 0.070 243.495 ;
    END
  END w_mask_in[1729]
  PIN w_mask_in[1730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.565 0.070 243.635 ;
    END
  END w_mask_in[1730]
  PIN w_mask_in[1731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.705 0.070 243.775 ;
    END
  END w_mask_in[1731]
  PIN w_mask_in[1732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.845 0.070 243.915 ;
    END
  END w_mask_in[1732]
  PIN w_mask_in[1733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 243.985 0.070 244.055 ;
    END
  END w_mask_in[1733]
  PIN w_mask_in[1734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.125 0.070 244.195 ;
    END
  END w_mask_in[1734]
  PIN w_mask_in[1735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.265 0.070 244.335 ;
    END
  END w_mask_in[1735]
  PIN w_mask_in[1736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.405 0.070 244.475 ;
    END
  END w_mask_in[1736]
  PIN w_mask_in[1737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.545 0.070 244.615 ;
    END
  END w_mask_in[1737]
  PIN w_mask_in[1738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.685 0.070 244.755 ;
    END
  END w_mask_in[1738]
  PIN w_mask_in[1739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.825 0.070 244.895 ;
    END
  END w_mask_in[1739]
  PIN w_mask_in[1740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.965 0.070 245.035 ;
    END
  END w_mask_in[1740]
  PIN w_mask_in[1741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.105 0.070 245.175 ;
    END
  END w_mask_in[1741]
  PIN w_mask_in[1742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.245 0.070 245.315 ;
    END
  END w_mask_in[1742]
  PIN w_mask_in[1743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.385 0.070 245.455 ;
    END
  END w_mask_in[1743]
  PIN w_mask_in[1744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.525 0.070 245.595 ;
    END
  END w_mask_in[1744]
  PIN w_mask_in[1745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.665 0.070 245.735 ;
    END
  END w_mask_in[1745]
  PIN w_mask_in[1746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.805 0.070 245.875 ;
    END
  END w_mask_in[1746]
  PIN w_mask_in[1747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 245.945 0.070 246.015 ;
    END
  END w_mask_in[1747]
  PIN w_mask_in[1748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.085 0.070 246.155 ;
    END
  END w_mask_in[1748]
  PIN w_mask_in[1749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.225 0.070 246.295 ;
    END
  END w_mask_in[1749]
  PIN w_mask_in[1750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.365 0.070 246.435 ;
    END
  END w_mask_in[1750]
  PIN w_mask_in[1751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.505 0.070 246.575 ;
    END
  END w_mask_in[1751]
  PIN w_mask_in[1752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.645 0.070 246.715 ;
    END
  END w_mask_in[1752]
  PIN w_mask_in[1753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.785 0.070 246.855 ;
    END
  END w_mask_in[1753]
  PIN w_mask_in[1754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.925 0.070 246.995 ;
    END
  END w_mask_in[1754]
  PIN w_mask_in[1755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.065 0.070 247.135 ;
    END
  END w_mask_in[1755]
  PIN w_mask_in[1756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.205 0.070 247.275 ;
    END
  END w_mask_in[1756]
  PIN w_mask_in[1757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.345 0.070 247.415 ;
    END
  END w_mask_in[1757]
  PIN w_mask_in[1758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.485 0.070 247.555 ;
    END
  END w_mask_in[1758]
  PIN w_mask_in[1759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.625 0.070 247.695 ;
    END
  END w_mask_in[1759]
  PIN w_mask_in[1760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.765 0.070 247.835 ;
    END
  END w_mask_in[1760]
  PIN w_mask_in[1761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.905 0.070 247.975 ;
    END
  END w_mask_in[1761]
  PIN w_mask_in[1762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.045 0.070 248.115 ;
    END
  END w_mask_in[1762]
  PIN w_mask_in[1763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.185 0.070 248.255 ;
    END
  END w_mask_in[1763]
  PIN w_mask_in[1764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.325 0.070 248.395 ;
    END
  END w_mask_in[1764]
  PIN w_mask_in[1765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.465 0.070 248.535 ;
    END
  END w_mask_in[1765]
  PIN w_mask_in[1766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.605 0.070 248.675 ;
    END
  END w_mask_in[1766]
  PIN w_mask_in[1767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.745 0.070 248.815 ;
    END
  END w_mask_in[1767]
  PIN w_mask_in[1768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 248.885 0.070 248.955 ;
    END
  END w_mask_in[1768]
  PIN w_mask_in[1769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.025 0.070 249.095 ;
    END
  END w_mask_in[1769]
  PIN w_mask_in[1770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.165 0.070 249.235 ;
    END
  END w_mask_in[1770]
  PIN w_mask_in[1771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.305 0.070 249.375 ;
    END
  END w_mask_in[1771]
  PIN w_mask_in[1772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.445 0.070 249.515 ;
    END
  END w_mask_in[1772]
  PIN w_mask_in[1773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.585 0.070 249.655 ;
    END
  END w_mask_in[1773]
  PIN w_mask_in[1774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.725 0.070 249.795 ;
    END
  END w_mask_in[1774]
  PIN w_mask_in[1775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.865 0.070 249.935 ;
    END
  END w_mask_in[1775]
  PIN w_mask_in[1776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.005 0.070 250.075 ;
    END
  END w_mask_in[1776]
  PIN w_mask_in[1777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.145 0.070 250.215 ;
    END
  END w_mask_in[1777]
  PIN w_mask_in[1778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.285 0.070 250.355 ;
    END
  END w_mask_in[1778]
  PIN w_mask_in[1779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.425 0.070 250.495 ;
    END
  END w_mask_in[1779]
  PIN w_mask_in[1780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.565 0.070 250.635 ;
    END
  END w_mask_in[1780]
  PIN w_mask_in[1781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.705 0.070 250.775 ;
    END
  END w_mask_in[1781]
  PIN w_mask_in[1782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.845 0.070 250.915 ;
    END
  END w_mask_in[1782]
  PIN w_mask_in[1783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.985 0.070 251.055 ;
    END
  END w_mask_in[1783]
  PIN w_mask_in[1784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.125 0.070 251.195 ;
    END
  END w_mask_in[1784]
  PIN w_mask_in[1785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.265 0.070 251.335 ;
    END
  END w_mask_in[1785]
  PIN w_mask_in[1786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.405 0.070 251.475 ;
    END
  END w_mask_in[1786]
  PIN w_mask_in[1787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.545 0.070 251.615 ;
    END
  END w_mask_in[1787]
  PIN w_mask_in[1788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.685 0.070 251.755 ;
    END
  END w_mask_in[1788]
  PIN w_mask_in[1789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.825 0.070 251.895 ;
    END
  END w_mask_in[1789]
  PIN w_mask_in[1790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.965 0.070 252.035 ;
    END
  END w_mask_in[1790]
  PIN w_mask_in[1791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.105 0.070 252.175 ;
    END
  END w_mask_in[1791]
  PIN w_mask_in[1792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.245 0.070 252.315 ;
    END
  END w_mask_in[1792]
  PIN w_mask_in[1793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.385 0.070 252.455 ;
    END
  END w_mask_in[1793]
  PIN w_mask_in[1794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.525 0.070 252.595 ;
    END
  END w_mask_in[1794]
  PIN w_mask_in[1795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.665 0.070 252.735 ;
    END
  END w_mask_in[1795]
  PIN w_mask_in[1796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.805 0.070 252.875 ;
    END
  END w_mask_in[1796]
  PIN w_mask_in[1797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.945 0.070 253.015 ;
    END
  END w_mask_in[1797]
  PIN w_mask_in[1798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.085 0.070 253.155 ;
    END
  END w_mask_in[1798]
  PIN w_mask_in[1799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.225 0.070 253.295 ;
    END
  END w_mask_in[1799]
  PIN w_mask_in[1800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.365 0.070 253.435 ;
    END
  END w_mask_in[1800]
  PIN w_mask_in[1801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.505 0.070 253.575 ;
    END
  END w_mask_in[1801]
  PIN w_mask_in[1802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.645 0.070 253.715 ;
    END
  END w_mask_in[1802]
  PIN w_mask_in[1803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.785 0.070 253.855 ;
    END
  END w_mask_in[1803]
  PIN w_mask_in[1804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.925 0.070 253.995 ;
    END
  END w_mask_in[1804]
  PIN w_mask_in[1805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.065 0.070 254.135 ;
    END
  END w_mask_in[1805]
  PIN w_mask_in[1806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.205 0.070 254.275 ;
    END
  END w_mask_in[1806]
  PIN w_mask_in[1807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.345 0.070 254.415 ;
    END
  END w_mask_in[1807]
  PIN w_mask_in[1808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.485 0.070 254.555 ;
    END
  END w_mask_in[1808]
  PIN w_mask_in[1809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.625 0.070 254.695 ;
    END
  END w_mask_in[1809]
  PIN w_mask_in[1810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.765 0.070 254.835 ;
    END
  END w_mask_in[1810]
  PIN w_mask_in[1811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.905 0.070 254.975 ;
    END
  END w_mask_in[1811]
  PIN w_mask_in[1812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.045 0.070 255.115 ;
    END
  END w_mask_in[1812]
  PIN w_mask_in[1813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.185 0.070 255.255 ;
    END
  END w_mask_in[1813]
  PIN w_mask_in[1814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.325 0.070 255.395 ;
    END
  END w_mask_in[1814]
  PIN w_mask_in[1815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.465 0.070 255.535 ;
    END
  END w_mask_in[1815]
  PIN w_mask_in[1816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.605 0.070 255.675 ;
    END
  END w_mask_in[1816]
  PIN w_mask_in[1817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.745 0.070 255.815 ;
    END
  END w_mask_in[1817]
  PIN w_mask_in[1818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.885 0.070 255.955 ;
    END
  END w_mask_in[1818]
  PIN w_mask_in[1819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.025 0.070 256.095 ;
    END
  END w_mask_in[1819]
  PIN w_mask_in[1820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.165 0.070 256.235 ;
    END
  END w_mask_in[1820]
  PIN w_mask_in[1821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.305 0.070 256.375 ;
    END
  END w_mask_in[1821]
  PIN w_mask_in[1822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.445 0.070 256.515 ;
    END
  END w_mask_in[1822]
  PIN w_mask_in[1823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.585 0.070 256.655 ;
    END
  END w_mask_in[1823]
  PIN w_mask_in[1824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.725 0.070 256.795 ;
    END
  END w_mask_in[1824]
  PIN w_mask_in[1825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.865 0.070 256.935 ;
    END
  END w_mask_in[1825]
  PIN w_mask_in[1826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.005 0.070 257.075 ;
    END
  END w_mask_in[1826]
  PIN w_mask_in[1827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.145 0.070 257.215 ;
    END
  END w_mask_in[1827]
  PIN w_mask_in[1828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.285 0.070 257.355 ;
    END
  END w_mask_in[1828]
  PIN w_mask_in[1829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.425 0.070 257.495 ;
    END
  END w_mask_in[1829]
  PIN w_mask_in[1830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.565 0.070 257.635 ;
    END
  END w_mask_in[1830]
  PIN w_mask_in[1831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.705 0.070 257.775 ;
    END
  END w_mask_in[1831]
  PIN w_mask_in[1832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.845 0.070 257.915 ;
    END
  END w_mask_in[1832]
  PIN w_mask_in[1833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.985 0.070 258.055 ;
    END
  END w_mask_in[1833]
  PIN w_mask_in[1834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.125 0.070 258.195 ;
    END
  END w_mask_in[1834]
  PIN w_mask_in[1835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.265 0.070 258.335 ;
    END
  END w_mask_in[1835]
  PIN w_mask_in[1836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.405 0.070 258.475 ;
    END
  END w_mask_in[1836]
  PIN w_mask_in[1837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.545 0.070 258.615 ;
    END
  END w_mask_in[1837]
  PIN w_mask_in[1838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.685 0.070 258.755 ;
    END
  END w_mask_in[1838]
  PIN w_mask_in[1839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.825 0.070 258.895 ;
    END
  END w_mask_in[1839]
  PIN w_mask_in[1840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.965 0.070 259.035 ;
    END
  END w_mask_in[1840]
  PIN w_mask_in[1841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.105 0.070 259.175 ;
    END
  END w_mask_in[1841]
  PIN w_mask_in[1842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.245 0.070 259.315 ;
    END
  END w_mask_in[1842]
  PIN w_mask_in[1843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.385 0.070 259.455 ;
    END
  END w_mask_in[1843]
  PIN w_mask_in[1844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.525 0.070 259.595 ;
    END
  END w_mask_in[1844]
  PIN w_mask_in[1845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.665 0.070 259.735 ;
    END
  END w_mask_in[1845]
  PIN w_mask_in[1846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.805 0.070 259.875 ;
    END
  END w_mask_in[1846]
  PIN w_mask_in[1847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.945 0.070 260.015 ;
    END
  END w_mask_in[1847]
  PIN w_mask_in[1848]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.085 0.070 260.155 ;
    END
  END w_mask_in[1848]
  PIN w_mask_in[1849]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.225 0.070 260.295 ;
    END
  END w_mask_in[1849]
  PIN w_mask_in[1850]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.365 0.070 260.435 ;
    END
  END w_mask_in[1850]
  PIN w_mask_in[1851]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.505 0.070 260.575 ;
    END
  END w_mask_in[1851]
  PIN w_mask_in[1852]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.645 0.070 260.715 ;
    END
  END w_mask_in[1852]
  PIN w_mask_in[1853]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.785 0.070 260.855 ;
    END
  END w_mask_in[1853]
  PIN w_mask_in[1854]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.925 0.070 260.995 ;
    END
  END w_mask_in[1854]
  PIN w_mask_in[1855]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.065 0.070 261.135 ;
    END
  END w_mask_in[1855]
  PIN w_mask_in[1856]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.205 0.070 261.275 ;
    END
  END w_mask_in[1856]
  PIN w_mask_in[1857]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.345 0.070 261.415 ;
    END
  END w_mask_in[1857]
  PIN w_mask_in[1858]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.485 0.070 261.555 ;
    END
  END w_mask_in[1858]
  PIN w_mask_in[1859]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.625 0.070 261.695 ;
    END
  END w_mask_in[1859]
  PIN w_mask_in[1860]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.765 0.070 261.835 ;
    END
  END w_mask_in[1860]
  PIN w_mask_in[1861]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 261.905 0.070 261.975 ;
    END
  END w_mask_in[1861]
  PIN w_mask_in[1862]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.045 0.070 262.115 ;
    END
  END w_mask_in[1862]
  PIN w_mask_in[1863]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.185 0.070 262.255 ;
    END
  END w_mask_in[1863]
  PIN w_mask_in[1864]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.325 0.070 262.395 ;
    END
  END w_mask_in[1864]
  PIN w_mask_in[1865]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.465 0.070 262.535 ;
    END
  END w_mask_in[1865]
  PIN w_mask_in[1866]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.605 0.070 262.675 ;
    END
  END w_mask_in[1866]
  PIN w_mask_in[1867]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.745 0.070 262.815 ;
    END
  END w_mask_in[1867]
  PIN w_mask_in[1868]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.885 0.070 262.955 ;
    END
  END w_mask_in[1868]
  PIN w_mask_in[1869]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.025 0.070 263.095 ;
    END
  END w_mask_in[1869]
  PIN w_mask_in[1870]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.165 0.070 263.235 ;
    END
  END w_mask_in[1870]
  PIN w_mask_in[1871]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.305 0.070 263.375 ;
    END
  END w_mask_in[1871]
  PIN w_mask_in[1872]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.445 0.070 263.515 ;
    END
  END w_mask_in[1872]
  PIN w_mask_in[1873]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.585 0.070 263.655 ;
    END
  END w_mask_in[1873]
  PIN w_mask_in[1874]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.725 0.070 263.795 ;
    END
  END w_mask_in[1874]
  PIN w_mask_in[1875]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.865 0.070 263.935 ;
    END
  END w_mask_in[1875]
  PIN w_mask_in[1876]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.005 0.070 264.075 ;
    END
  END w_mask_in[1876]
  PIN w_mask_in[1877]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.145 0.070 264.215 ;
    END
  END w_mask_in[1877]
  PIN w_mask_in[1878]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.285 0.070 264.355 ;
    END
  END w_mask_in[1878]
  PIN w_mask_in[1879]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.425 0.070 264.495 ;
    END
  END w_mask_in[1879]
  PIN w_mask_in[1880]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.565 0.070 264.635 ;
    END
  END w_mask_in[1880]
  PIN w_mask_in[1881]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.705 0.070 264.775 ;
    END
  END w_mask_in[1881]
  PIN w_mask_in[1882]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.845 0.070 264.915 ;
    END
  END w_mask_in[1882]
  PIN w_mask_in[1883]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.985 0.070 265.055 ;
    END
  END w_mask_in[1883]
  PIN w_mask_in[1884]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.125 0.070 265.195 ;
    END
  END w_mask_in[1884]
  PIN w_mask_in[1885]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.265 0.070 265.335 ;
    END
  END w_mask_in[1885]
  PIN w_mask_in[1886]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.405 0.070 265.475 ;
    END
  END w_mask_in[1886]
  PIN w_mask_in[1887]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.545 0.070 265.615 ;
    END
  END w_mask_in[1887]
  PIN w_mask_in[1888]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.685 0.070 265.755 ;
    END
  END w_mask_in[1888]
  PIN w_mask_in[1889]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.825 0.070 265.895 ;
    END
  END w_mask_in[1889]
  PIN w_mask_in[1890]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 265.965 0.070 266.035 ;
    END
  END w_mask_in[1890]
  PIN w_mask_in[1891]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.105 0.070 266.175 ;
    END
  END w_mask_in[1891]
  PIN w_mask_in[1892]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.245 0.070 266.315 ;
    END
  END w_mask_in[1892]
  PIN w_mask_in[1893]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.385 0.070 266.455 ;
    END
  END w_mask_in[1893]
  PIN w_mask_in[1894]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.525 0.070 266.595 ;
    END
  END w_mask_in[1894]
  PIN w_mask_in[1895]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.665 0.070 266.735 ;
    END
  END w_mask_in[1895]
  PIN w_mask_in[1896]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.805 0.070 266.875 ;
    END
  END w_mask_in[1896]
  PIN w_mask_in[1897]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.945 0.070 267.015 ;
    END
  END w_mask_in[1897]
  PIN w_mask_in[1898]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.085 0.070 267.155 ;
    END
  END w_mask_in[1898]
  PIN w_mask_in[1899]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.225 0.070 267.295 ;
    END
  END w_mask_in[1899]
  PIN w_mask_in[1900]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.365 0.070 267.435 ;
    END
  END w_mask_in[1900]
  PIN w_mask_in[1901]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.505 0.070 267.575 ;
    END
  END w_mask_in[1901]
  PIN w_mask_in[1902]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.645 0.070 267.715 ;
    END
  END w_mask_in[1902]
  PIN w_mask_in[1903]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.785 0.070 267.855 ;
    END
  END w_mask_in[1903]
  PIN w_mask_in[1904]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.925 0.070 267.995 ;
    END
  END w_mask_in[1904]
  PIN w_mask_in[1905]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.065 0.070 268.135 ;
    END
  END w_mask_in[1905]
  PIN w_mask_in[1906]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.205 0.070 268.275 ;
    END
  END w_mask_in[1906]
  PIN w_mask_in[1907]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.345 0.070 268.415 ;
    END
  END w_mask_in[1907]
  PIN w_mask_in[1908]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.485 0.070 268.555 ;
    END
  END w_mask_in[1908]
  PIN w_mask_in[1909]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.625 0.070 268.695 ;
    END
  END w_mask_in[1909]
  PIN w_mask_in[1910]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.765 0.070 268.835 ;
    END
  END w_mask_in[1910]
  PIN w_mask_in[1911]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.905 0.070 268.975 ;
    END
  END w_mask_in[1911]
  PIN w_mask_in[1912]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.045 0.070 269.115 ;
    END
  END w_mask_in[1912]
  PIN w_mask_in[1913]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.185 0.070 269.255 ;
    END
  END w_mask_in[1913]
  PIN w_mask_in[1914]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.325 0.070 269.395 ;
    END
  END w_mask_in[1914]
  PIN w_mask_in[1915]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.465 0.070 269.535 ;
    END
  END w_mask_in[1915]
  PIN w_mask_in[1916]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.605 0.070 269.675 ;
    END
  END w_mask_in[1916]
  PIN w_mask_in[1917]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.745 0.070 269.815 ;
    END
  END w_mask_in[1917]
  PIN w_mask_in[1918]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.885 0.070 269.955 ;
    END
  END w_mask_in[1918]
  PIN w_mask_in[1919]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.025 0.070 270.095 ;
    END
  END w_mask_in[1919]
  PIN w_mask_in[1920]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.165 0.070 270.235 ;
    END
  END w_mask_in[1920]
  PIN w_mask_in[1921]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.305 0.070 270.375 ;
    END
  END w_mask_in[1921]
  PIN w_mask_in[1922]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.445 0.070 270.515 ;
    END
  END w_mask_in[1922]
  PIN w_mask_in[1923]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.585 0.070 270.655 ;
    END
  END w_mask_in[1923]
  PIN w_mask_in[1924]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.725 0.070 270.795 ;
    END
  END w_mask_in[1924]
  PIN w_mask_in[1925]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.865 0.070 270.935 ;
    END
  END w_mask_in[1925]
  PIN w_mask_in[1926]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.005 0.070 271.075 ;
    END
  END w_mask_in[1926]
  PIN w_mask_in[1927]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.145 0.070 271.215 ;
    END
  END w_mask_in[1927]
  PIN w_mask_in[1928]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.285 0.070 271.355 ;
    END
  END w_mask_in[1928]
  PIN w_mask_in[1929]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.425 0.070 271.495 ;
    END
  END w_mask_in[1929]
  PIN w_mask_in[1930]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.565 0.070 271.635 ;
    END
  END w_mask_in[1930]
  PIN w_mask_in[1931]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.705 0.070 271.775 ;
    END
  END w_mask_in[1931]
  PIN w_mask_in[1932]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.845 0.070 271.915 ;
    END
  END w_mask_in[1932]
  PIN w_mask_in[1933]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.985 0.070 272.055 ;
    END
  END w_mask_in[1933]
  PIN w_mask_in[1934]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.125 0.070 272.195 ;
    END
  END w_mask_in[1934]
  PIN w_mask_in[1935]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.265 0.070 272.335 ;
    END
  END w_mask_in[1935]
  PIN w_mask_in[1936]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.405 0.070 272.475 ;
    END
  END w_mask_in[1936]
  PIN w_mask_in[1937]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.545 0.070 272.615 ;
    END
  END w_mask_in[1937]
  PIN w_mask_in[1938]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.685 0.070 272.755 ;
    END
  END w_mask_in[1938]
  PIN w_mask_in[1939]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.825 0.070 272.895 ;
    END
  END w_mask_in[1939]
  PIN w_mask_in[1940]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.965 0.070 273.035 ;
    END
  END w_mask_in[1940]
  PIN w_mask_in[1941]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.105 0.070 273.175 ;
    END
  END w_mask_in[1941]
  PIN w_mask_in[1942]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.245 0.070 273.315 ;
    END
  END w_mask_in[1942]
  PIN w_mask_in[1943]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.385 0.070 273.455 ;
    END
  END w_mask_in[1943]
  PIN w_mask_in[1944]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.525 0.070 273.595 ;
    END
  END w_mask_in[1944]
  PIN w_mask_in[1945]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.665 0.070 273.735 ;
    END
  END w_mask_in[1945]
  PIN w_mask_in[1946]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.805 0.070 273.875 ;
    END
  END w_mask_in[1946]
  PIN w_mask_in[1947]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.945 0.070 274.015 ;
    END
  END w_mask_in[1947]
  PIN w_mask_in[1948]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.085 0.070 274.155 ;
    END
  END w_mask_in[1948]
  PIN w_mask_in[1949]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.225 0.070 274.295 ;
    END
  END w_mask_in[1949]
  PIN w_mask_in[1950]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.365 0.070 274.435 ;
    END
  END w_mask_in[1950]
  PIN w_mask_in[1951]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.505 0.070 274.575 ;
    END
  END w_mask_in[1951]
  PIN w_mask_in[1952]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.645 0.070 274.715 ;
    END
  END w_mask_in[1952]
  PIN w_mask_in[1953]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.785 0.070 274.855 ;
    END
  END w_mask_in[1953]
  PIN w_mask_in[1954]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.925 0.070 274.995 ;
    END
  END w_mask_in[1954]
  PIN w_mask_in[1955]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.065 0.070 275.135 ;
    END
  END w_mask_in[1955]
  PIN w_mask_in[1956]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.205 0.070 275.275 ;
    END
  END w_mask_in[1956]
  PIN w_mask_in[1957]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.345 0.070 275.415 ;
    END
  END w_mask_in[1957]
  PIN w_mask_in[1958]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.485 0.070 275.555 ;
    END
  END w_mask_in[1958]
  PIN w_mask_in[1959]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.625 0.070 275.695 ;
    END
  END w_mask_in[1959]
  PIN w_mask_in[1960]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.765 0.070 275.835 ;
    END
  END w_mask_in[1960]
  PIN w_mask_in[1961]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 275.905 0.070 275.975 ;
    END
  END w_mask_in[1961]
  PIN w_mask_in[1962]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.045 0.070 276.115 ;
    END
  END w_mask_in[1962]
  PIN w_mask_in[1963]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.185 0.070 276.255 ;
    END
  END w_mask_in[1963]
  PIN w_mask_in[1964]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.325 0.070 276.395 ;
    END
  END w_mask_in[1964]
  PIN w_mask_in[1965]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.465 0.070 276.535 ;
    END
  END w_mask_in[1965]
  PIN w_mask_in[1966]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.605 0.070 276.675 ;
    END
  END w_mask_in[1966]
  PIN w_mask_in[1967]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.745 0.070 276.815 ;
    END
  END w_mask_in[1967]
  PIN w_mask_in[1968]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.885 0.070 276.955 ;
    END
  END w_mask_in[1968]
  PIN w_mask_in[1969]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.025 0.070 277.095 ;
    END
  END w_mask_in[1969]
  PIN w_mask_in[1970]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.165 0.070 277.235 ;
    END
  END w_mask_in[1970]
  PIN w_mask_in[1971]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.305 0.070 277.375 ;
    END
  END w_mask_in[1971]
  PIN w_mask_in[1972]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.445 0.070 277.515 ;
    END
  END w_mask_in[1972]
  PIN w_mask_in[1973]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.585 0.070 277.655 ;
    END
  END w_mask_in[1973]
  PIN w_mask_in[1974]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.725 0.070 277.795 ;
    END
  END w_mask_in[1974]
  PIN w_mask_in[1975]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.865 0.070 277.935 ;
    END
  END w_mask_in[1975]
  PIN w_mask_in[1976]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.005 0.070 278.075 ;
    END
  END w_mask_in[1976]
  PIN w_mask_in[1977]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.145 0.070 278.215 ;
    END
  END w_mask_in[1977]
  PIN w_mask_in[1978]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.285 0.070 278.355 ;
    END
  END w_mask_in[1978]
  PIN w_mask_in[1979]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.425 0.070 278.495 ;
    END
  END w_mask_in[1979]
  PIN w_mask_in[1980]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.565 0.070 278.635 ;
    END
  END w_mask_in[1980]
  PIN w_mask_in[1981]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.705 0.070 278.775 ;
    END
  END w_mask_in[1981]
  PIN w_mask_in[1982]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.845 0.070 278.915 ;
    END
  END w_mask_in[1982]
  PIN w_mask_in[1983]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 278.985 0.070 279.055 ;
    END
  END w_mask_in[1983]
  PIN w_mask_in[1984]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.125 0.070 279.195 ;
    END
  END w_mask_in[1984]
  PIN w_mask_in[1985]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.265 0.070 279.335 ;
    END
  END w_mask_in[1985]
  PIN w_mask_in[1986]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.405 0.070 279.475 ;
    END
  END w_mask_in[1986]
  PIN w_mask_in[1987]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.545 0.070 279.615 ;
    END
  END w_mask_in[1987]
  PIN w_mask_in[1988]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.685 0.070 279.755 ;
    END
  END w_mask_in[1988]
  PIN w_mask_in[1989]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.825 0.070 279.895 ;
    END
  END w_mask_in[1989]
  PIN w_mask_in[1990]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.965 0.070 280.035 ;
    END
  END w_mask_in[1990]
  PIN w_mask_in[1991]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.105 0.070 280.175 ;
    END
  END w_mask_in[1991]
  PIN w_mask_in[1992]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.245 0.070 280.315 ;
    END
  END w_mask_in[1992]
  PIN w_mask_in[1993]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.385 0.070 280.455 ;
    END
  END w_mask_in[1993]
  PIN w_mask_in[1994]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.525 0.070 280.595 ;
    END
  END w_mask_in[1994]
  PIN w_mask_in[1995]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.665 0.070 280.735 ;
    END
  END w_mask_in[1995]
  PIN w_mask_in[1996]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.805 0.070 280.875 ;
    END
  END w_mask_in[1996]
  PIN w_mask_in[1997]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.945 0.070 281.015 ;
    END
  END w_mask_in[1997]
  PIN w_mask_in[1998]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.085 0.070 281.155 ;
    END
  END w_mask_in[1998]
  PIN w_mask_in[1999]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.225 0.070 281.295 ;
    END
  END w_mask_in[1999]
  PIN w_mask_in[2000]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.365 0.070 281.435 ;
    END
  END w_mask_in[2000]
  PIN w_mask_in[2001]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.505 0.070 281.575 ;
    END
  END w_mask_in[2001]
  PIN w_mask_in[2002]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.645 0.070 281.715 ;
    END
  END w_mask_in[2002]
  PIN w_mask_in[2003]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.785 0.070 281.855 ;
    END
  END w_mask_in[2003]
  PIN w_mask_in[2004]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 281.925 0.070 281.995 ;
    END
  END w_mask_in[2004]
  PIN w_mask_in[2005]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.065 0.070 282.135 ;
    END
  END w_mask_in[2005]
  PIN w_mask_in[2006]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.205 0.070 282.275 ;
    END
  END w_mask_in[2006]
  PIN w_mask_in[2007]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.345 0.070 282.415 ;
    END
  END w_mask_in[2007]
  PIN w_mask_in[2008]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.485 0.070 282.555 ;
    END
  END w_mask_in[2008]
  PIN w_mask_in[2009]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.625 0.070 282.695 ;
    END
  END w_mask_in[2009]
  PIN w_mask_in[2010]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.765 0.070 282.835 ;
    END
  END w_mask_in[2010]
  PIN w_mask_in[2011]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.905 0.070 282.975 ;
    END
  END w_mask_in[2011]
  PIN w_mask_in[2012]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.045 0.070 283.115 ;
    END
  END w_mask_in[2012]
  PIN w_mask_in[2013]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.185 0.070 283.255 ;
    END
  END w_mask_in[2013]
  PIN w_mask_in[2014]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.325 0.070 283.395 ;
    END
  END w_mask_in[2014]
  PIN w_mask_in[2015]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.465 0.070 283.535 ;
    END
  END w_mask_in[2015]
  PIN w_mask_in[2016]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.605 0.070 283.675 ;
    END
  END w_mask_in[2016]
  PIN w_mask_in[2017]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.745 0.070 283.815 ;
    END
  END w_mask_in[2017]
  PIN w_mask_in[2018]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 283.885 0.070 283.955 ;
    END
  END w_mask_in[2018]
  PIN w_mask_in[2019]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.025 0.070 284.095 ;
    END
  END w_mask_in[2019]
  PIN w_mask_in[2020]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.165 0.070 284.235 ;
    END
  END w_mask_in[2020]
  PIN w_mask_in[2021]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.305 0.070 284.375 ;
    END
  END w_mask_in[2021]
  PIN w_mask_in[2022]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.445 0.070 284.515 ;
    END
  END w_mask_in[2022]
  PIN w_mask_in[2023]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.585 0.070 284.655 ;
    END
  END w_mask_in[2023]
  PIN w_mask_in[2024]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.725 0.070 284.795 ;
    END
  END w_mask_in[2024]
  PIN w_mask_in[2025]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.865 0.070 284.935 ;
    END
  END w_mask_in[2025]
  PIN w_mask_in[2026]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.005 0.070 285.075 ;
    END
  END w_mask_in[2026]
  PIN w_mask_in[2027]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.145 0.070 285.215 ;
    END
  END w_mask_in[2027]
  PIN w_mask_in[2028]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.285 0.070 285.355 ;
    END
  END w_mask_in[2028]
  PIN w_mask_in[2029]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.425 0.070 285.495 ;
    END
  END w_mask_in[2029]
  PIN w_mask_in[2030]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.565 0.070 285.635 ;
    END
  END w_mask_in[2030]
  PIN w_mask_in[2031]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.705 0.070 285.775 ;
    END
  END w_mask_in[2031]
  PIN w_mask_in[2032]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.845 0.070 285.915 ;
    END
  END w_mask_in[2032]
  PIN w_mask_in[2033]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.985 0.070 286.055 ;
    END
  END w_mask_in[2033]
  PIN w_mask_in[2034]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.125 0.070 286.195 ;
    END
  END w_mask_in[2034]
  PIN w_mask_in[2035]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.265 0.070 286.335 ;
    END
  END w_mask_in[2035]
  PIN w_mask_in[2036]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.405 0.070 286.475 ;
    END
  END w_mask_in[2036]
  PIN w_mask_in[2037]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.545 0.070 286.615 ;
    END
  END w_mask_in[2037]
  PIN w_mask_in[2038]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.685 0.070 286.755 ;
    END
  END w_mask_in[2038]
  PIN w_mask_in[2039]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.825 0.070 286.895 ;
    END
  END w_mask_in[2039]
  PIN w_mask_in[2040]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 286.965 0.070 287.035 ;
    END
  END w_mask_in[2040]
  PIN w_mask_in[2041]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.105 0.070 287.175 ;
    END
  END w_mask_in[2041]
  PIN w_mask_in[2042]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.245 0.070 287.315 ;
    END
  END w_mask_in[2042]
  PIN w_mask_in[2043]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.385 0.070 287.455 ;
    END
  END w_mask_in[2043]
  PIN w_mask_in[2044]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.525 0.070 287.595 ;
    END
  END w_mask_in[2044]
  PIN w_mask_in[2045]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.665 0.070 287.735 ;
    END
  END w_mask_in[2045]
  PIN w_mask_in[2046]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.805 0.070 287.875 ;
    END
  END w_mask_in[2046]
  PIN w_mask_in[2047]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.945 0.070 288.015 ;
    END
  END w_mask_in[2047]
  PIN w_mask_in[2048]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.085 0.070 288.155 ;
    END
  END w_mask_in[2048]
  PIN w_mask_in[2049]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.225 0.070 288.295 ;
    END
  END w_mask_in[2049]
  PIN w_mask_in[2050]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.365 0.070 288.435 ;
    END
  END w_mask_in[2050]
  PIN w_mask_in[2051]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.505 0.070 288.575 ;
    END
  END w_mask_in[2051]
  PIN w_mask_in[2052]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.645 0.070 288.715 ;
    END
  END w_mask_in[2052]
  PIN w_mask_in[2053]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.785 0.070 288.855 ;
    END
  END w_mask_in[2053]
  PIN w_mask_in[2054]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.925 0.070 288.995 ;
    END
  END w_mask_in[2054]
  PIN w_mask_in[2055]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.065 0.070 289.135 ;
    END
  END w_mask_in[2055]
  PIN w_mask_in[2056]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.205 0.070 289.275 ;
    END
  END w_mask_in[2056]
  PIN w_mask_in[2057]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.345 0.070 289.415 ;
    END
  END w_mask_in[2057]
  PIN w_mask_in[2058]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.485 0.070 289.555 ;
    END
  END w_mask_in[2058]
  PIN w_mask_in[2059]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.625 0.070 289.695 ;
    END
  END w_mask_in[2059]
  PIN w_mask_in[2060]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.765 0.070 289.835 ;
    END
  END w_mask_in[2060]
  PIN w_mask_in[2061]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.905 0.070 289.975 ;
    END
  END w_mask_in[2061]
  PIN w_mask_in[2062]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.045 0.070 290.115 ;
    END
  END w_mask_in[2062]
  PIN w_mask_in[2063]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.185 0.070 290.255 ;
    END
  END w_mask_in[2063]
  PIN w_mask_in[2064]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.325 0.070 290.395 ;
    END
  END w_mask_in[2064]
  PIN w_mask_in[2065]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.465 0.070 290.535 ;
    END
  END w_mask_in[2065]
  PIN w_mask_in[2066]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.605 0.070 290.675 ;
    END
  END w_mask_in[2066]
  PIN w_mask_in[2067]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.745 0.070 290.815 ;
    END
  END w_mask_in[2067]
  PIN w_mask_in[2068]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 290.885 0.070 290.955 ;
    END
  END w_mask_in[2068]
  PIN w_mask_in[2069]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.025 0.070 291.095 ;
    END
  END w_mask_in[2069]
  PIN w_mask_in[2070]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.165 0.070 291.235 ;
    END
  END w_mask_in[2070]
  PIN w_mask_in[2071]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.305 0.070 291.375 ;
    END
  END w_mask_in[2071]
  PIN w_mask_in[2072]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.445 0.070 291.515 ;
    END
  END w_mask_in[2072]
  PIN w_mask_in[2073]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.585 0.070 291.655 ;
    END
  END w_mask_in[2073]
  PIN w_mask_in[2074]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.725 0.070 291.795 ;
    END
  END w_mask_in[2074]
  PIN w_mask_in[2075]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.865 0.070 291.935 ;
    END
  END w_mask_in[2075]
  PIN w_mask_in[2076]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.005 0.070 292.075 ;
    END
  END w_mask_in[2076]
  PIN w_mask_in[2077]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.145 0.070 292.215 ;
    END
  END w_mask_in[2077]
  PIN w_mask_in[2078]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.285 0.070 292.355 ;
    END
  END w_mask_in[2078]
  PIN w_mask_in[2079]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.425 0.070 292.495 ;
    END
  END w_mask_in[2079]
  PIN w_mask_in[2080]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.565 0.070 292.635 ;
    END
  END w_mask_in[2080]
  PIN w_mask_in[2081]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.705 0.070 292.775 ;
    END
  END w_mask_in[2081]
  PIN w_mask_in[2082]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.845 0.070 292.915 ;
    END
  END w_mask_in[2082]
  PIN w_mask_in[2083]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.985 0.070 293.055 ;
    END
  END w_mask_in[2083]
  PIN w_mask_in[2084]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.125 0.070 293.195 ;
    END
  END w_mask_in[2084]
  PIN w_mask_in[2085]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.265 0.070 293.335 ;
    END
  END w_mask_in[2085]
  PIN w_mask_in[2086]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.405 0.070 293.475 ;
    END
  END w_mask_in[2086]
  PIN w_mask_in[2087]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.545 0.070 293.615 ;
    END
  END w_mask_in[2087]
  PIN w_mask_in[2088]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.685 0.070 293.755 ;
    END
  END w_mask_in[2088]
  PIN w_mask_in[2089]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.825 0.070 293.895 ;
    END
  END w_mask_in[2089]
  PIN w_mask_in[2090]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 293.965 0.070 294.035 ;
    END
  END w_mask_in[2090]
  PIN w_mask_in[2091]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.105 0.070 294.175 ;
    END
  END w_mask_in[2091]
  PIN w_mask_in[2092]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.245 0.070 294.315 ;
    END
  END w_mask_in[2092]
  PIN w_mask_in[2093]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.385 0.070 294.455 ;
    END
  END w_mask_in[2093]
  PIN w_mask_in[2094]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.525 0.070 294.595 ;
    END
  END w_mask_in[2094]
  PIN w_mask_in[2095]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.665 0.070 294.735 ;
    END
  END w_mask_in[2095]
  PIN w_mask_in[2096]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.805 0.070 294.875 ;
    END
  END w_mask_in[2096]
  PIN w_mask_in[2097]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.945 0.070 295.015 ;
    END
  END w_mask_in[2097]
  PIN w_mask_in[2098]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.085 0.070 295.155 ;
    END
  END w_mask_in[2098]
  PIN w_mask_in[2099]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.225 0.070 295.295 ;
    END
  END w_mask_in[2099]
  PIN w_mask_in[2100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.365 0.070 295.435 ;
    END
  END w_mask_in[2100]
  PIN w_mask_in[2101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.505 0.070 295.575 ;
    END
  END w_mask_in[2101]
  PIN w_mask_in[2102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.645 0.070 295.715 ;
    END
  END w_mask_in[2102]
  PIN w_mask_in[2103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.785 0.070 295.855 ;
    END
  END w_mask_in[2103]
  PIN w_mask_in[2104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 295.925 0.070 295.995 ;
    END
  END w_mask_in[2104]
  PIN w_mask_in[2105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.065 0.070 296.135 ;
    END
  END w_mask_in[2105]
  PIN w_mask_in[2106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.205 0.070 296.275 ;
    END
  END w_mask_in[2106]
  PIN w_mask_in[2107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.345 0.070 296.415 ;
    END
  END w_mask_in[2107]
  PIN w_mask_in[2108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.485 0.070 296.555 ;
    END
  END w_mask_in[2108]
  PIN w_mask_in[2109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.625 0.070 296.695 ;
    END
  END w_mask_in[2109]
  PIN w_mask_in[2110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.765 0.070 296.835 ;
    END
  END w_mask_in[2110]
  PIN w_mask_in[2111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.905 0.070 296.975 ;
    END
  END w_mask_in[2111]
  PIN w_mask_in[2112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.045 0.070 297.115 ;
    END
  END w_mask_in[2112]
  PIN w_mask_in[2113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.185 0.070 297.255 ;
    END
  END w_mask_in[2113]
  PIN w_mask_in[2114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.325 0.070 297.395 ;
    END
  END w_mask_in[2114]
  PIN w_mask_in[2115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.465 0.070 297.535 ;
    END
  END w_mask_in[2115]
  PIN w_mask_in[2116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.605 0.070 297.675 ;
    END
  END w_mask_in[2116]
  PIN w_mask_in[2117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.745 0.070 297.815 ;
    END
  END w_mask_in[2117]
  PIN w_mask_in[2118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.885 0.070 297.955 ;
    END
  END w_mask_in[2118]
  PIN w_mask_in[2119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.025 0.070 298.095 ;
    END
  END w_mask_in[2119]
  PIN w_mask_in[2120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.165 0.070 298.235 ;
    END
  END w_mask_in[2120]
  PIN w_mask_in[2121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.305 0.070 298.375 ;
    END
  END w_mask_in[2121]
  PIN w_mask_in[2122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.445 0.070 298.515 ;
    END
  END w_mask_in[2122]
  PIN w_mask_in[2123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.585 0.070 298.655 ;
    END
  END w_mask_in[2123]
  PIN w_mask_in[2124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.725 0.070 298.795 ;
    END
  END w_mask_in[2124]
  PIN w_mask_in[2125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 298.865 0.070 298.935 ;
    END
  END w_mask_in[2125]
  PIN w_mask_in[2126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.005 0.070 299.075 ;
    END
  END w_mask_in[2126]
  PIN w_mask_in[2127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.145 0.070 299.215 ;
    END
  END w_mask_in[2127]
  PIN w_mask_in[2128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.285 0.070 299.355 ;
    END
  END w_mask_in[2128]
  PIN w_mask_in[2129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.425 0.070 299.495 ;
    END
  END w_mask_in[2129]
  PIN w_mask_in[2130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.565 0.070 299.635 ;
    END
  END w_mask_in[2130]
  PIN w_mask_in[2131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.705 0.070 299.775 ;
    END
  END w_mask_in[2131]
  PIN w_mask_in[2132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.845 0.070 299.915 ;
    END
  END w_mask_in[2132]
  PIN w_mask_in[2133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.985 0.070 300.055 ;
    END
  END w_mask_in[2133]
  PIN w_mask_in[2134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.125 0.070 300.195 ;
    END
  END w_mask_in[2134]
  PIN w_mask_in[2135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.265 0.070 300.335 ;
    END
  END w_mask_in[2135]
  PIN w_mask_in[2136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.405 0.070 300.475 ;
    END
  END w_mask_in[2136]
  PIN w_mask_in[2137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.545 0.070 300.615 ;
    END
  END w_mask_in[2137]
  PIN w_mask_in[2138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.685 0.070 300.755 ;
    END
  END w_mask_in[2138]
  PIN w_mask_in[2139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.825 0.070 300.895 ;
    END
  END w_mask_in[2139]
  PIN w_mask_in[2140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.965 0.070 301.035 ;
    END
  END w_mask_in[2140]
  PIN w_mask_in[2141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.105 0.070 301.175 ;
    END
  END w_mask_in[2141]
  PIN w_mask_in[2142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.245 0.070 301.315 ;
    END
  END w_mask_in[2142]
  PIN w_mask_in[2143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.385 0.070 301.455 ;
    END
  END w_mask_in[2143]
  PIN w_mask_in[2144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.525 0.070 301.595 ;
    END
  END w_mask_in[2144]
  PIN w_mask_in[2145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.665 0.070 301.735 ;
    END
  END w_mask_in[2145]
  PIN w_mask_in[2146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.805 0.070 301.875 ;
    END
  END w_mask_in[2146]
  PIN w_mask_in[2147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 301.945 0.070 302.015 ;
    END
  END w_mask_in[2147]
  PIN w_mask_in[2148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.085 0.070 302.155 ;
    END
  END w_mask_in[2148]
  PIN w_mask_in[2149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.225 0.070 302.295 ;
    END
  END w_mask_in[2149]
  PIN w_mask_in[2150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.365 0.070 302.435 ;
    END
  END w_mask_in[2150]
  PIN w_mask_in[2151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.505 0.070 302.575 ;
    END
  END w_mask_in[2151]
  PIN w_mask_in[2152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.645 0.070 302.715 ;
    END
  END w_mask_in[2152]
  PIN w_mask_in[2153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.785 0.070 302.855 ;
    END
  END w_mask_in[2153]
  PIN w_mask_in[2154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.925 0.070 302.995 ;
    END
  END w_mask_in[2154]
  PIN w_mask_in[2155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.065 0.070 303.135 ;
    END
  END w_mask_in[2155]
  PIN w_mask_in[2156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.205 0.070 303.275 ;
    END
  END w_mask_in[2156]
  PIN w_mask_in[2157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.345 0.070 303.415 ;
    END
  END w_mask_in[2157]
  PIN w_mask_in[2158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.485 0.070 303.555 ;
    END
  END w_mask_in[2158]
  PIN w_mask_in[2159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.625 0.070 303.695 ;
    END
  END w_mask_in[2159]
  PIN w_mask_in[2160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.765 0.070 303.835 ;
    END
  END w_mask_in[2160]
  PIN w_mask_in[2161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.905 0.070 303.975 ;
    END
  END w_mask_in[2161]
  PIN w_mask_in[2162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.045 0.070 304.115 ;
    END
  END w_mask_in[2162]
  PIN w_mask_in[2163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.185 0.070 304.255 ;
    END
  END w_mask_in[2163]
  PIN w_mask_in[2164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.325 0.070 304.395 ;
    END
  END w_mask_in[2164]
  PIN w_mask_in[2165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.465 0.070 304.535 ;
    END
  END w_mask_in[2165]
  PIN w_mask_in[2166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.605 0.070 304.675 ;
    END
  END w_mask_in[2166]
  PIN w_mask_in[2167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.745 0.070 304.815 ;
    END
  END w_mask_in[2167]
  PIN w_mask_in[2168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.885 0.070 304.955 ;
    END
  END w_mask_in[2168]
  PIN w_mask_in[2169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.025 0.070 305.095 ;
    END
  END w_mask_in[2169]
  PIN w_mask_in[2170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.165 0.070 305.235 ;
    END
  END w_mask_in[2170]
  PIN w_mask_in[2171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.305 0.070 305.375 ;
    END
  END w_mask_in[2171]
  PIN w_mask_in[2172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.445 0.070 305.515 ;
    END
  END w_mask_in[2172]
  PIN w_mask_in[2173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.585 0.070 305.655 ;
    END
  END w_mask_in[2173]
  PIN w_mask_in[2174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.725 0.070 305.795 ;
    END
  END w_mask_in[2174]
  PIN w_mask_in[2175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 305.865 0.070 305.935 ;
    END
  END w_mask_in[2175]
  PIN w_mask_in[2176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.005 0.070 306.075 ;
    END
  END w_mask_in[2176]
  PIN w_mask_in[2177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.145 0.070 306.215 ;
    END
  END w_mask_in[2177]
  PIN w_mask_in[2178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.285 0.070 306.355 ;
    END
  END w_mask_in[2178]
  PIN w_mask_in[2179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.425 0.070 306.495 ;
    END
  END w_mask_in[2179]
  PIN w_mask_in[2180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.565 0.070 306.635 ;
    END
  END w_mask_in[2180]
  PIN w_mask_in[2181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.705 0.070 306.775 ;
    END
  END w_mask_in[2181]
  PIN w_mask_in[2182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.845 0.070 306.915 ;
    END
  END w_mask_in[2182]
  PIN w_mask_in[2183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.985 0.070 307.055 ;
    END
  END w_mask_in[2183]
  PIN w_mask_in[2184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.125 0.070 307.195 ;
    END
  END w_mask_in[2184]
  PIN w_mask_in[2185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.265 0.070 307.335 ;
    END
  END w_mask_in[2185]
  PIN w_mask_in[2186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.405 0.070 307.475 ;
    END
  END w_mask_in[2186]
  PIN w_mask_in[2187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.545 0.070 307.615 ;
    END
  END w_mask_in[2187]
  PIN w_mask_in[2188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.685 0.070 307.755 ;
    END
  END w_mask_in[2188]
  PIN w_mask_in[2189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.825 0.070 307.895 ;
    END
  END w_mask_in[2189]
  PIN w_mask_in[2190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.965 0.070 308.035 ;
    END
  END w_mask_in[2190]
  PIN w_mask_in[2191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.105 0.070 308.175 ;
    END
  END w_mask_in[2191]
  PIN w_mask_in[2192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.245 0.070 308.315 ;
    END
  END w_mask_in[2192]
  PIN w_mask_in[2193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.385 0.070 308.455 ;
    END
  END w_mask_in[2193]
  PIN w_mask_in[2194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.525 0.070 308.595 ;
    END
  END w_mask_in[2194]
  PIN w_mask_in[2195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.665 0.070 308.735 ;
    END
  END w_mask_in[2195]
  PIN w_mask_in[2196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.805 0.070 308.875 ;
    END
  END w_mask_in[2196]
  PIN w_mask_in[2197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 308.945 0.070 309.015 ;
    END
  END w_mask_in[2197]
  PIN w_mask_in[2198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.085 0.070 309.155 ;
    END
  END w_mask_in[2198]
  PIN w_mask_in[2199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.225 0.070 309.295 ;
    END
  END w_mask_in[2199]
  PIN w_mask_in[2200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.365 0.070 309.435 ;
    END
  END w_mask_in[2200]
  PIN w_mask_in[2201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.505 0.070 309.575 ;
    END
  END w_mask_in[2201]
  PIN w_mask_in[2202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.645 0.070 309.715 ;
    END
  END w_mask_in[2202]
  PIN w_mask_in[2203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.785 0.070 309.855 ;
    END
  END w_mask_in[2203]
  PIN w_mask_in[2204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.925 0.070 309.995 ;
    END
  END w_mask_in[2204]
  PIN w_mask_in[2205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.065 0.070 310.135 ;
    END
  END w_mask_in[2205]
  PIN w_mask_in[2206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.205 0.070 310.275 ;
    END
  END w_mask_in[2206]
  PIN w_mask_in[2207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.345 0.070 310.415 ;
    END
  END w_mask_in[2207]
  PIN w_mask_in[2208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.485 0.070 310.555 ;
    END
  END w_mask_in[2208]
  PIN w_mask_in[2209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.625 0.070 310.695 ;
    END
  END w_mask_in[2209]
  PIN w_mask_in[2210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.765 0.070 310.835 ;
    END
  END w_mask_in[2210]
  PIN w_mask_in[2211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 310.905 0.070 310.975 ;
    END
  END w_mask_in[2211]
  PIN w_mask_in[2212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.045 0.070 311.115 ;
    END
  END w_mask_in[2212]
  PIN w_mask_in[2213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.185 0.070 311.255 ;
    END
  END w_mask_in[2213]
  PIN w_mask_in[2214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.325 0.070 311.395 ;
    END
  END w_mask_in[2214]
  PIN w_mask_in[2215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.465 0.070 311.535 ;
    END
  END w_mask_in[2215]
  PIN w_mask_in[2216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.605 0.070 311.675 ;
    END
  END w_mask_in[2216]
  PIN w_mask_in[2217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.745 0.070 311.815 ;
    END
  END w_mask_in[2217]
  PIN w_mask_in[2218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 311.885 0.070 311.955 ;
    END
  END w_mask_in[2218]
  PIN w_mask_in[2219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.025 0.070 312.095 ;
    END
  END w_mask_in[2219]
  PIN w_mask_in[2220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.165 0.070 312.235 ;
    END
  END w_mask_in[2220]
  PIN w_mask_in[2221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.305 0.070 312.375 ;
    END
  END w_mask_in[2221]
  PIN w_mask_in[2222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.445 0.070 312.515 ;
    END
  END w_mask_in[2222]
  PIN w_mask_in[2223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.585 0.070 312.655 ;
    END
  END w_mask_in[2223]
  PIN w_mask_in[2224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.725 0.070 312.795 ;
    END
  END w_mask_in[2224]
  PIN w_mask_in[2225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.865 0.070 312.935 ;
    END
  END w_mask_in[2225]
  PIN w_mask_in[2226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.005 0.070 313.075 ;
    END
  END w_mask_in[2226]
  PIN w_mask_in[2227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.145 0.070 313.215 ;
    END
  END w_mask_in[2227]
  PIN w_mask_in[2228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.285 0.070 313.355 ;
    END
  END w_mask_in[2228]
  PIN w_mask_in[2229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.425 0.070 313.495 ;
    END
  END w_mask_in[2229]
  PIN w_mask_in[2230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.565 0.070 313.635 ;
    END
  END w_mask_in[2230]
  PIN w_mask_in[2231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.705 0.070 313.775 ;
    END
  END w_mask_in[2231]
  PIN w_mask_in[2232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.845 0.070 313.915 ;
    END
  END w_mask_in[2232]
  PIN w_mask_in[2233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 313.985 0.070 314.055 ;
    END
  END w_mask_in[2233]
  PIN w_mask_in[2234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.125 0.070 314.195 ;
    END
  END w_mask_in[2234]
  PIN w_mask_in[2235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.265 0.070 314.335 ;
    END
  END w_mask_in[2235]
  PIN w_mask_in[2236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.405 0.070 314.475 ;
    END
  END w_mask_in[2236]
  PIN w_mask_in[2237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.545 0.070 314.615 ;
    END
  END w_mask_in[2237]
  PIN w_mask_in[2238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.685 0.070 314.755 ;
    END
  END w_mask_in[2238]
  PIN w_mask_in[2239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.825 0.070 314.895 ;
    END
  END w_mask_in[2239]
  PIN w_mask_in[2240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.965 0.070 315.035 ;
    END
  END w_mask_in[2240]
  PIN w_mask_in[2241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.105 0.070 315.175 ;
    END
  END w_mask_in[2241]
  PIN w_mask_in[2242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.245 0.070 315.315 ;
    END
  END w_mask_in[2242]
  PIN w_mask_in[2243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.385 0.070 315.455 ;
    END
  END w_mask_in[2243]
  PIN w_mask_in[2244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.525 0.070 315.595 ;
    END
  END w_mask_in[2244]
  PIN w_mask_in[2245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.665 0.070 315.735 ;
    END
  END w_mask_in[2245]
  PIN w_mask_in[2246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.805 0.070 315.875 ;
    END
  END w_mask_in[2246]
  PIN w_mask_in[2247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 315.945 0.070 316.015 ;
    END
  END w_mask_in[2247]
  PIN w_mask_in[2248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.085 0.070 316.155 ;
    END
  END w_mask_in[2248]
  PIN w_mask_in[2249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.225 0.070 316.295 ;
    END
  END w_mask_in[2249]
  PIN w_mask_in[2250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.365 0.070 316.435 ;
    END
  END w_mask_in[2250]
  PIN w_mask_in[2251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.505 0.070 316.575 ;
    END
  END w_mask_in[2251]
  PIN w_mask_in[2252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.645 0.070 316.715 ;
    END
  END w_mask_in[2252]
  PIN w_mask_in[2253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.785 0.070 316.855 ;
    END
  END w_mask_in[2253]
  PIN w_mask_in[2254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 316.925 0.070 316.995 ;
    END
  END w_mask_in[2254]
  PIN w_mask_in[2255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.065 0.070 317.135 ;
    END
  END w_mask_in[2255]
  PIN w_mask_in[2256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.205 0.070 317.275 ;
    END
  END w_mask_in[2256]
  PIN w_mask_in[2257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.345 0.070 317.415 ;
    END
  END w_mask_in[2257]
  PIN w_mask_in[2258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.485 0.070 317.555 ;
    END
  END w_mask_in[2258]
  PIN w_mask_in[2259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.625 0.070 317.695 ;
    END
  END w_mask_in[2259]
  PIN w_mask_in[2260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.765 0.070 317.835 ;
    END
  END w_mask_in[2260]
  PIN w_mask_in[2261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.905 0.070 317.975 ;
    END
  END w_mask_in[2261]
  PIN w_mask_in[2262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.045 0.070 318.115 ;
    END
  END w_mask_in[2262]
  PIN w_mask_in[2263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.185 0.070 318.255 ;
    END
  END w_mask_in[2263]
  PIN w_mask_in[2264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.325 0.070 318.395 ;
    END
  END w_mask_in[2264]
  PIN w_mask_in[2265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.465 0.070 318.535 ;
    END
  END w_mask_in[2265]
  PIN w_mask_in[2266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.605 0.070 318.675 ;
    END
  END w_mask_in[2266]
  PIN w_mask_in[2267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.745 0.070 318.815 ;
    END
  END w_mask_in[2267]
  PIN w_mask_in[2268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 318.885 0.070 318.955 ;
    END
  END w_mask_in[2268]
  PIN w_mask_in[2269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.025 0.070 319.095 ;
    END
  END w_mask_in[2269]
  PIN w_mask_in[2270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.165 0.070 319.235 ;
    END
  END w_mask_in[2270]
  PIN w_mask_in[2271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.305 0.070 319.375 ;
    END
  END w_mask_in[2271]
  PIN w_mask_in[2272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.445 0.070 319.515 ;
    END
  END w_mask_in[2272]
  PIN w_mask_in[2273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.585 0.070 319.655 ;
    END
  END w_mask_in[2273]
  PIN w_mask_in[2274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.725 0.070 319.795 ;
    END
  END w_mask_in[2274]
  PIN w_mask_in[2275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 319.865 0.070 319.935 ;
    END
  END w_mask_in[2275]
  PIN w_mask_in[2276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.005 0.070 320.075 ;
    END
  END w_mask_in[2276]
  PIN w_mask_in[2277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.145 0.070 320.215 ;
    END
  END w_mask_in[2277]
  PIN w_mask_in[2278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.285 0.070 320.355 ;
    END
  END w_mask_in[2278]
  PIN w_mask_in[2279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.425 0.070 320.495 ;
    END
  END w_mask_in[2279]
  PIN w_mask_in[2280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.565 0.070 320.635 ;
    END
  END w_mask_in[2280]
  PIN w_mask_in[2281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.705 0.070 320.775 ;
    END
  END w_mask_in[2281]
  PIN w_mask_in[2282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.845 0.070 320.915 ;
    END
  END w_mask_in[2282]
  PIN w_mask_in[2283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.985 0.070 321.055 ;
    END
  END w_mask_in[2283]
  PIN w_mask_in[2284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.125 0.070 321.195 ;
    END
  END w_mask_in[2284]
  PIN w_mask_in[2285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.265 0.070 321.335 ;
    END
  END w_mask_in[2285]
  PIN w_mask_in[2286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.405 0.070 321.475 ;
    END
  END w_mask_in[2286]
  PIN w_mask_in[2287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.545 0.070 321.615 ;
    END
  END w_mask_in[2287]
  PIN w_mask_in[2288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.685 0.070 321.755 ;
    END
  END w_mask_in[2288]
  PIN w_mask_in[2289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.825 0.070 321.895 ;
    END
  END w_mask_in[2289]
  PIN w_mask_in[2290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 321.965 0.070 322.035 ;
    END
  END w_mask_in[2290]
  PIN w_mask_in[2291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.105 0.070 322.175 ;
    END
  END w_mask_in[2291]
  PIN w_mask_in[2292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.245 0.070 322.315 ;
    END
  END w_mask_in[2292]
  PIN w_mask_in[2293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.385 0.070 322.455 ;
    END
  END w_mask_in[2293]
  PIN w_mask_in[2294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.525 0.070 322.595 ;
    END
  END w_mask_in[2294]
  PIN w_mask_in[2295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.665 0.070 322.735 ;
    END
  END w_mask_in[2295]
  PIN w_mask_in[2296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.805 0.070 322.875 ;
    END
  END w_mask_in[2296]
  PIN w_mask_in[2297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.945 0.070 323.015 ;
    END
  END w_mask_in[2297]
  PIN w_mask_in[2298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.085 0.070 323.155 ;
    END
  END w_mask_in[2298]
  PIN w_mask_in[2299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.225 0.070 323.295 ;
    END
  END w_mask_in[2299]
  PIN w_mask_in[2300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.365 0.070 323.435 ;
    END
  END w_mask_in[2300]
  PIN w_mask_in[2301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.505 0.070 323.575 ;
    END
  END w_mask_in[2301]
  PIN w_mask_in[2302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.645 0.070 323.715 ;
    END
  END w_mask_in[2302]
  PIN w_mask_in[2303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.785 0.070 323.855 ;
    END
  END w_mask_in[2303]
  PIN w_mask_in[2304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.925 0.070 323.995 ;
    END
  END w_mask_in[2304]
  PIN w_mask_in[2305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.065 0.070 324.135 ;
    END
  END w_mask_in[2305]
  PIN w_mask_in[2306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.205 0.070 324.275 ;
    END
  END w_mask_in[2306]
  PIN w_mask_in[2307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.345 0.070 324.415 ;
    END
  END w_mask_in[2307]
  PIN w_mask_in[2308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.485 0.070 324.555 ;
    END
  END w_mask_in[2308]
  PIN w_mask_in[2309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.625 0.070 324.695 ;
    END
  END w_mask_in[2309]
  PIN w_mask_in[2310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.765 0.070 324.835 ;
    END
  END w_mask_in[2310]
  PIN w_mask_in[2311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 324.905 0.070 324.975 ;
    END
  END w_mask_in[2311]
  PIN w_mask_in[2312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.045 0.070 325.115 ;
    END
  END w_mask_in[2312]
  PIN w_mask_in[2313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.185 0.070 325.255 ;
    END
  END w_mask_in[2313]
  PIN w_mask_in[2314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.325 0.070 325.395 ;
    END
  END w_mask_in[2314]
  PIN w_mask_in[2315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.465 0.070 325.535 ;
    END
  END w_mask_in[2315]
  PIN w_mask_in[2316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.605 0.070 325.675 ;
    END
  END w_mask_in[2316]
  PIN w_mask_in[2317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.745 0.070 325.815 ;
    END
  END w_mask_in[2317]
  PIN w_mask_in[2318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.885 0.070 325.955 ;
    END
  END w_mask_in[2318]
  PIN w_mask_in[2319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.025 0.070 326.095 ;
    END
  END w_mask_in[2319]
  PIN w_mask_in[2320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.165 0.070 326.235 ;
    END
  END w_mask_in[2320]
  PIN w_mask_in[2321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.305 0.070 326.375 ;
    END
  END w_mask_in[2321]
  PIN w_mask_in[2322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.445 0.070 326.515 ;
    END
  END w_mask_in[2322]
  PIN w_mask_in[2323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.585 0.070 326.655 ;
    END
  END w_mask_in[2323]
  PIN w_mask_in[2324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.725 0.070 326.795 ;
    END
  END w_mask_in[2324]
  PIN w_mask_in[2325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.865 0.070 326.935 ;
    END
  END w_mask_in[2325]
  PIN w_mask_in[2326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.005 0.070 327.075 ;
    END
  END w_mask_in[2326]
  PIN w_mask_in[2327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.145 0.070 327.215 ;
    END
  END w_mask_in[2327]
  PIN w_mask_in[2328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.285 0.070 327.355 ;
    END
  END w_mask_in[2328]
  PIN w_mask_in[2329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.425 0.070 327.495 ;
    END
  END w_mask_in[2329]
  PIN w_mask_in[2330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.565 0.070 327.635 ;
    END
  END w_mask_in[2330]
  PIN w_mask_in[2331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.705 0.070 327.775 ;
    END
  END w_mask_in[2331]
  PIN w_mask_in[2332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.845 0.070 327.915 ;
    END
  END w_mask_in[2332]
  PIN w_mask_in[2333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 327.985 0.070 328.055 ;
    END
  END w_mask_in[2333]
  PIN w_mask_in[2334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.125 0.070 328.195 ;
    END
  END w_mask_in[2334]
  PIN w_mask_in[2335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.265 0.070 328.335 ;
    END
  END w_mask_in[2335]
  PIN w_mask_in[2336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.405 0.070 328.475 ;
    END
  END w_mask_in[2336]
  PIN w_mask_in[2337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.545 0.070 328.615 ;
    END
  END w_mask_in[2337]
  PIN w_mask_in[2338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.685 0.070 328.755 ;
    END
  END w_mask_in[2338]
  PIN w_mask_in[2339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.825 0.070 328.895 ;
    END
  END w_mask_in[2339]
  PIN w_mask_in[2340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 328.965 0.070 329.035 ;
    END
  END w_mask_in[2340]
  PIN w_mask_in[2341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.105 0.070 329.175 ;
    END
  END w_mask_in[2341]
  PIN w_mask_in[2342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.245 0.070 329.315 ;
    END
  END w_mask_in[2342]
  PIN w_mask_in[2343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.385 0.070 329.455 ;
    END
  END w_mask_in[2343]
  PIN w_mask_in[2344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.525 0.070 329.595 ;
    END
  END w_mask_in[2344]
  PIN w_mask_in[2345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.665 0.070 329.735 ;
    END
  END w_mask_in[2345]
  PIN w_mask_in[2346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.805 0.070 329.875 ;
    END
  END w_mask_in[2346]
  PIN w_mask_in[2347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.945 0.070 330.015 ;
    END
  END w_mask_in[2347]
  PIN w_mask_in[2348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.085 0.070 330.155 ;
    END
  END w_mask_in[2348]
  PIN w_mask_in[2349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.225 0.070 330.295 ;
    END
  END w_mask_in[2349]
  PIN w_mask_in[2350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.365 0.070 330.435 ;
    END
  END w_mask_in[2350]
  PIN w_mask_in[2351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.505 0.070 330.575 ;
    END
  END w_mask_in[2351]
  PIN w_mask_in[2352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.645 0.070 330.715 ;
    END
  END w_mask_in[2352]
  PIN w_mask_in[2353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.785 0.070 330.855 ;
    END
  END w_mask_in[2353]
  PIN w_mask_in[2354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 330.925 0.070 330.995 ;
    END
  END w_mask_in[2354]
  PIN w_mask_in[2355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.065 0.070 331.135 ;
    END
  END w_mask_in[2355]
  PIN w_mask_in[2356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.205 0.070 331.275 ;
    END
  END w_mask_in[2356]
  PIN w_mask_in[2357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.345 0.070 331.415 ;
    END
  END w_mask_in[2357]
  PIN w_mask_in[2358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.485 0.070 331.555 ;
    END
  END w_mask_in[2358]
  PIN w_mask_in[2359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.625 0.070 331.695 ;
    END
  END w_mask_in[2359]
  PIN w_mask_in[2360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.765 0.070 331.835 ;
    END
  END w_mask_in[2360]
  PIN w_mask_in[2361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.905 0.070 331.975 ;
    END
  END w_mask_in[2361]
  PIN w_mask_in[2362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.045 0.070 332.115 ;
    END
  END w_mask_in[2362]
  PIN w_mask_in[2363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.185 0.070 332.255 ;
    END
  END w_mask_in[2363]
  PIN w_mask_in[2364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.325 0.070 332.395 ;
    END
  END w_mask_in[2364]
  PIN w_mask_in[2365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.465 0.070 332.535 ;
    END
  END w_mask_in[2365]
  PIN w_mask_in[2366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.605 0.070 332.675 ;
    END
  END w_mask_in[2366]
  PIN w_mask_in[2367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.745 0.070 332.815 ;
    END
  END w_mask_in[2367]
  PIN w_mask_in[2368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.885 0.070 332.955 ;
    END
  END w_mask_in[2368]
  PIN w_mask_in[2369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.025 0.070 333.095 ;
    END
  END w_mask_in[2369]
  PIN w_mask_in[2370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.165 0.070 333.235 ;
    END
  END w_mask_in[2370]
  PIN w_mask_in[2371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.305 0.070 333.375 ;
    END
  END w_mask_in[2371]
  PIN w_mask_in[2372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.445 0.070 333.515 ;
    END
  END w_mask_in[2372]
  PIN w_mask_in[2373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.585 0.070 333.655 ;
    END
  END w_mask_in[2373]
  PIN w_mask_in[2374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.725 0.070 333.795 ;
    END
  END w_mask_in[2374]
  PIN w_mask_in[2375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.865 0.070 333.935 ;
    END
  END w_mask_in[2375]
  PIN w_mask_in[2376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.005 0.070 334.075 ;
    END
  END w_mask_in[2376]
  PIN w_mask_in[2377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.145 0.070 334.215 ;
    END
  END w_mask_in[2377]
  PIN w_mask_in[2378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.285 0.070 334.355 ;
    END
  END w_mask_in[2378]
  PIN w_mask_in[2379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.425 0.070 334.495 ;
    END
  END w_mask_in[2379]
  PIN w_mask_in[2380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.565 0.070 334.635 ;
    END
  END w_mask_in[2380]
  PIN w_mask_in[2381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.705 0.070 334.775 ;
    END
  END w_mask_in[2381]
  PIN w_mask_in[2382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.845 0.070 334.915 ;
    END
  END w_mask_in[2382]
  PIN w_mask_in[2383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 334.985 0.070 335.055 ;
    END
  END w_mask_in[2383]
  PIN w_mask_in[2384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.125 0.070 335.195 ;
    END
  END w_mask_in[2384]
  PIN w_mask_in[2385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.265 0.070 335.335 ;
    END
  END w_mask_in[2385]
  PIN w_mask_in[2386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.405 0.070 335.475 ;
    END
  END w_mask_in[2386]
  PIN w_mask_in[2387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.545 0.070 335.615 ;
    END
  END w_mask_in[2387]
  PIN w_mask_in[2388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.685 0.070 335.755 ;
    END
  END w_mask_in[2388]
  PIN w_mask_in[2389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.825 0.070 335.895 ;
    END
  END w_mask_in[2389]
  PIN w_mask_in[2390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.965 0.070 336.035 ;
    END
  END w_mask_in[2390]
  PIN w_mask_in[2391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.105 0.070 336.175 ;
    END
  END w_mask_in[2391]
  PIN w_mask_in[2392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.245 0.070 336.315 ;
    END
  END w_mask_in[2392]
  PIN w_mask_in[2393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.385 0.070 336.455 ;
    END
  END w_mask_in[2393]
  PIN w_mask_in[2394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.525 0.070 336.595 ;
    END
  END w_mask_in[2394]
  PIN w_mask_in[2395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.665 0.070 336.735 ;
    END
  END w_mask_in[2395]
  PIN w_mask_in[2396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.805 0.070 336.875 ;
    END
  END w_mask_in[2396]
  PIN w_mask_in[2397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.945 0.070 337.015 ;
    END
  END w_mask_in[2397]
  PIN w_mask_in[2398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.085 0.070 337.155 ;
    END
  END w_mask_in[2398]
  PIN w_mask_in[2399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.225 0.070 337.295 ;
    END
  END w_mask_in[2399]
  PIN w_mask_in[2400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.365 0.070 337.435 ;
    END
  END w_mask_in[2400]
  PIN w_mask_in[2401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.505 0.070 337.575 ;
    END
  END w_mask_in[2401]
  PIN w_mask_in[2402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.645 0.070 337.715 ;
    END
  END w_mask_in[2402]
  PIN w_mask_in[2403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.785 0.070 337.855 ;
    END
  END w_mask_in[2403]
  PIN w_mask_in[2404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 337.925 0.070 337.995 ;
    END
  END w_mask_in[2404]
  PIN w_mask_in[2405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.065 0.070 338.135 ;
    END
  END w_mask_in[2405]
  PIN w_mask_in[2406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.205 0.070 338.275 ;
    END
  END w_mask_in[2406]
  PIN w_mask_in[2407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.345 0.070 338.415 ;
    END
  END w_mask_in[2407]
  PIN w_mask_in[2408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.485 0.070 338.555 ;
    END
  END w_mask_in[2408]
  PIN w_mask_in[2409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.625 0.070 338.695 ;
    END
  END w_mask_in[2409]
  PIN w_mask_in[2410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.765 0.070 338.835 ;
    END
  END w_mask_in[2410]
  PIN w_mask_in[2411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.905 0.070 338.975 ;
    END
  END w_mask_in[2411]
  PIN w_mask_in[2412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.045 0.070 339.115 ;
    END
  END w_mask_in[2412]
  PIN w_mask_in[2413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.185 0.070 339.255 ;
    END
  END w_mask_in[2413]
  PIN w_mask_in[2414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.325 0.070 339.395 ;
    END
  END w_mask_in[2414]
  PIN w_mask_in[2415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.465 0.070 339.535 ;
    END
  END w_mask_in[2415]
  PIN w_mask_in[2416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.605 0.070 339.675 ;
    END
  END w_mask_in[2416]
  PIN w_mask_in[2417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.745 0.070 339.815 ;
    END
  END w_mask_in[2417]
  PIN w_mask_in[2418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 339.885 0.070 339.955 ;
    END
  END w_mask_in[2418]
  PIN w_mask_in[2419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.025 0.070 340.095 ;
    END
  END w_mask_in[2419]
  PIN w_mask_in[2420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.165 0.070 340.235 ;
    END
  END w_mask_in[2420]
  PIN w_mask_in[2421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.305 0.070 340.375 ;
    END
  END w_mask_in[2421]
  PIN w_mask_in[2422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.445 0.070 340.515 ;
    END
  END w_mask_in[2422]
  PIN w_mask_in[2423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.585 0.070 340.655 ;
    END
  END w_mask_in[2423]
  PIN w_mask_in[2424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.725 0.070 340.795 ;
    END
  END w_mask_in[2424]
  PIN w_mask_in[2425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 340.865 0.070 340.935 ;
    END
  END w_mask_in[2425]
  PIN w_mask_in[2426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.005 0.070 341.075 ;
    END
  END w_mask_in[2426]
  PIN w_mask_in[2427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.145 0.070 341.215 ;
    END
  END w_mask_in[2427]
  PIN w_mask_in[2428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.285 0.070 341.355 ;
    END
  END w_mask_in[2428]
  PIN w_mask_in[2429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.425 0.070 341.495 ;
    END
  END w_mask_in[2429]
  PIN w_mask_in[2430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.565 0.070 341.635 ;
    END
  END w_mask_in[2430]
  PIN w_mask_in[2431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.705 0.070 341.775 ;
    END
  END w_mask_in[2431]
  PIN w_mask_in[2432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.845 0.070 341.915 ;
    END
  END w_mask_in[2432]
  PIN w_mask_in[2433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.985 0.070 342.055 ;
    END
  END w_mask_in[2433]
  PIN w_mask_in[2434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.125 0.070 342.195 ;
    END
  END w_mask_in[2434]
  PIN w_mask_in[2435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.265 0.070 342.335 ;
    END
  END w_mask_in[2435]
  PIN w_mask_in[2436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.405 0.070 342.475 ;
    END
  END w_mask_in[2436]
  PIN w_mask_in[2437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.545 0.070 342.615 ;
    END
  END w_mask_in[2437]
  PIN w_mask_in[2438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.685 0.070 342.755 ;
    END
  END w_mask_in[2438]
  PIN w_mask_in[2439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.825 0.070 342.895 ;
    END
  END w_mask_in[2439]
  PIN w_mask_in[2440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 342.965 0.070 343.035 ;
    END
  END w_mask_in[2440]
  PIN w_mask_in[2441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.105 0.070 343.175 ;
    END
  END w_mask_in[2441]
  PIN w_mask_in[2442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.245 0.070 343.315 ;
    END
  END w_mask_in[2442]
  PIN w_mask_in[2443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.385 0.070 343.455 ;
    END
  END w_mask_in[2443]
  PIN w_mask_in[2444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.525 0.070 343.595 ;
    END
  END w_mask_in[2444]
  PIN w_mask_in[2445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.665 0.070 343.735 ;
    END
  END w_mask_in[2445]
  PIN w_mask_in[2446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.805 0.070 343.875 ;
    END
  END w_mask_in[2446]
  PIN w_mask_in[2447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.945 0.070 344.015 ;
    END
  END w_mask_in[2447]
  PIN w_mask_in[2448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.085 0.070 344.155 ;
    END
  END w_mask_in[2448]
  PIN w_mask_in[2449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.225 0.070 344.295 ;
    END
  END w_mask_in[2449]
  PIN w_mask_in[2450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.365 0.070 344.435 ;
    END
  END w_mask_in[2450]
  PIN w_mask_in[2451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.505 0.070 344.575 ;
    END
  END w_mask_in[2451]
  PIN w_mask_in[2452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.645 0.070 344.715 ;
    END
  END w_mask_in[2452]
  PIN w_mask_in[2453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.785 0.070 344.855 ;
    END
  END w_mask_in[2453]
  PIN w_mask_in[2454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.925 0.070 344.995 ;
    END
  END w_mask_in[2454]
  PIN w_mask_in[2455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.065 0.070 345.135 ;
    END
  END w_mask_in[2455]
  PIN w_mask_in[2456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.205 0.070 345.275 ;
    END
  END w_mask_in[2456]
  PIN w_mask_in[2457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.345 0.070 345.415 ;
    END
  END w_mask_in[2457]
  PIN w_mask_in[2458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.485 0.070 345.555 ;
    END
  END w_mask_in[2458]
  PIN w_mask_in[2459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.625 0.070 345.695 ;
    END
  END w_mask_in[2459]
  PIN w_mask_in[2460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.765 0.070 345.835 ;
    END
  END w_mask_in[2460]
  PIN w_mask_in[2461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 345.905 0.070 345.975 ;
    END
  END w_mask_in[2461]
  PIN w_mask_in[2462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.045 0.070 346.115 ;
    END
  END w_mask_in[2462]
  PIN w_mask_in[2463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.185 0.070 346.255 ;
    END
  END w_mask_in[2463]
  PIN w_mask_in[2464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.325 0.070 346.395 ;
    END
  END w_mask_in[2464]
  PIN w_mask_in[2465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.465 0.070 346.535 ;
    END
  END w_mask_in[2465]
  PIN w_mask_in[2466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.605 0.070 346.675 ;
    END
  END w_mask_in[2466]
  PIN w_mask_in[2467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.745 0.070 346.815 ;
    END
  END w_mask_in[2467]
  PIN w_mask_in[2468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.885 0.070 346.955 ;
    END
  END w_mask_in[2468]
  PIN w_mask_in[2469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.025 0.070 347.095 ;
    END
  END w_mask_in[2469]
  PIN w_mask_in[2470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.165 0.070 347.235 ;
    END
  END w_mask_in[2470]
  PIN w_mask_in[2471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.305 0.070 347.375 ;
    END
  END w_mask_in[2471]
  PIN w_mask_in[2472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.445 0.070 347.515 ;
    END
  END w_mask_in[2472]
  PIN w_mask_in[2473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.585 0.070 347.655 ;
    END
  END w_mask_in[2473]
  PIN w_mask_in[2474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.725 0.070 347.795 ;
    END
  END w_mask_in[2474]
  PIN w_mask_in[2475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.865 0.070 347.935 ;
    END
  END w_mask_in[2475]
  PIN w_mask_in[2476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.005 0.070 348.075 ;
    END
  END w_mask_in[2476]
  PIN w_mask_in[2477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.145 0.070 348.215 ;
    END
  END w_mask_in[2477]
  PIN w_mask_in[2478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.285 0.070 348.355 ;
    END
  END w_mask_in[2478]
  PIN w_mask_in[2479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.425 0.070 348.495 ;
    END
  END w_mask_in[2479]
  PIN w_mask_in[2480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.565 0.070 348.635 ;
    END
  END w_mask_in[2480]
  PIN w_mask_in[2481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.705 0.070 348.775 ;
    END
  END w_mask_in[2481]
  PIN w_mask_in[2482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.845 0.070 348.915 ;
    END
  END w_mask_in[2482]
  PIN w_mask_in[2483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.985 0.070 349.055 ;
    END
  END w_mask_in[2483]
  PIN w_mask_in[2484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.125 0.070 349.195 ;
    END
  END w_mask_in[2484]
  PIN w_mask_in[2485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.265 0.070 349.335 ;
    END
  END w_mask_in[2485]
  PIN w_mask_in[2486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.405 0.070 349.475 ;
    END
  END w_mask_in[2486]
  PIN w_mask_in[2487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.545 0.070 349.615 ;
    END
  END w_mask_in[2487]
  PIN w_mask_in[2488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.685 0.070 349.755 ;
    END
  END w_mask_in[2488]
  PIN w_mask_in[2489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.825 0.070 349.895 ;
    END
  END w_mask_in[2489]
  PIN w_mask_in[2490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 349.965 0.070 350.035 ;
    END
  END w_mask_in[2490]
  PIN w_mask_in[2491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.105 0.070 350.175 ;
    END
  END w_mask_in[2491]
  PIN w_mask_in[2492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.245 0.070 350.315 ;
    END
  END w_mask_in[2492]
  PIN w_mask_in[2493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.385 0.070 350.455 ;
    END
  END w_mask_in[2493]
  PIN w_mask_in[2494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.525 0.070 350.595 ;
    END
  END w_mask_in[2494]
  PIN w_mask_in[2495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.665 0.070 350.735 ;
    END
  END w_mask_in[2495]
  PIN w_mask_in[2496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.805 0.070 350.875 ;
    END
  END w_mask_in[2496]
  PIN w_mask_in[2497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.945 0.070 351.015 ;
    END
  END w_mask_in[2497]
  PIN w_mask_in[2498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.085 0.070 351.155 ;
    END
  END w_mask_in[2498]
  PIN w_mask_in[2499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.225 0.070 351.295 ;
    END
  END w_mask_in[2499]
  PIN w_mask_in[2500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.365 0.070 351.435 ;
    END
  END w_mask_in[2500]
  PIN w_mask_in[2501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.505 0.070 351.575 ;
    END
  END w_mask_in[2501]
  PIN w_mask_in[2502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.645 0.070 351.715 ;
    END
  END w_mask_in[2502]
  PIN w_mask_in[2503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.785 0.070 351.855 ;
    END
  END w_mask_in[2503]
  PIN w_mask_in[2504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.925 0.070 351.995 ;
    END
  END w_mask_in[2504]
  PIN w_mask_in[2505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.065 0.070 352.135 ;
    END
  END w_mask_in[2505]
  PIN w_mask_in[2506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.205 0.070 352.275 ;
    END
  END w_mask_in[2506]
  PIN w_mask_in[2507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.345 0.070 352.415 ;
    END
  END w_mask_in[2507]
  PIN w_mask_in[2508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.485 0.070 352.555 ;
    END
  END w_mask_in[2508]
  PIN w_mask_in[2509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.625 0.070 352.695 ;
    END
  END w_mask_in[2509]
  PIN w_mask_in[2510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.765 0.070 352.835 ;
    END
  END w_mask_in[2510]
  PIN w_mask_in[2511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 352.905 0.070 352.975 ;
    END
  END w_mask_in[2511]
  PIN w_mask_in[2512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.045 0.070 353.115 ;
    END
  END w_mask_in[2512]
  PIN w_mask_in[2513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.185 0.070 353.255 ;
    END
  END w_mask_in[2513]
  PIN w_mask_in[2514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.325 0.070 353.395 ;
    END
  END w_mask_in[2514]
  PIN w_mask_in[2515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.465 0.070 353.535 ;
    END
  END w_mask_in[2515]
  PIN w_mask_in[2516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.605 0.070 353.675 ;
    END
  END w_mask_in[2516]
  PIN w_mask_in[2517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.745 0.070 353.815 ;
    END
  END w_mask_in[2517]
  PIN w_mask_in[2518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.885 0.070 353.955 ;
    END
  END w_mask_in[2518]
  PIN w_mask_in[2519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.025 0.070 354.095 ;
    END
  END w_mask_in[2519]
  PIN w_mask_in[2520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.165 0.070 354.235 ;
    END
  END w_mask_in[2520]
  PIN w_mask_in[2521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.305 0.070 354.375 ;
    END
  END w_mask_in[2521]
  PIN w_mask_in[2522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.445 0.070 354.515 ;
    END
  END w_mask_in[2522]
  PIN w_mask_in[2523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.585 0.070 354.655 ;
    END
  END w_mask_in[2523]
  PIN w_mask_in[2524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.725 0.070 354.795 ;
    END
  END w_mask_in[2524]
  PIN w_mask_in[2525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 354.865 0.070 354.935 ;
    END
  END w_mask_in[2525]
  PIN w_mask_in[2526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.005 0.070 355.075 ;
    END
  END w_mask_in[2526]
  PIN w_mask_in[2527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.145 0.070 355.215 ;
    END
  END w_mask_in[2527]
  PIN w_mask_in[2528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.285 0.070 355.355 ;
    END
  END w_mask_in[2528]
  PIN w_mask_in[2529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.425 0.070 355.495 ;
    END
  END w_mask_in[2529]
  PIN w_mask_in[2530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.565 0.070 355.635 ;
    END
  END w_mask_in[2530]
  PIN w_mask_in[2531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.705 0.070 355.775 ;
    END
  END w_mask_in[2531]
  PIN w_mask_in[2532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.845 0.070 355.915 ;
    END
  END w_mask_in[2532]
  PIN w_mask_in[2533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 355.985 0.070 356.055 ;
    END
  END w_mask_in[2533]
  PIN w_mask_in[2534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.125 0.070 356.195 ;
    END
  END w_mask_in[2534]
  PIN w_mask_in[2535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.265 0.070 356.335 ;
    END
  END w_mask_in[2535]
  PIN w_mask_in[2536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.405 0.070 356.475 ;
    END
  END w_mask_in[2536]
  PIN w_mask_in[2537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.545 0.070 356.615 ;
    END
  END w_mask_in[2537]
  PIN w_mask_in[2538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.685 0.070 356.755 ;
    END
  END w_mask_in[2538]
  PIN w_mask_in[2539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.825 0.070 356.895 ;
    END
  END w_mask_in[2539]
  PIN w_mask_in[2540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.965 0.070 357.035 ;
    END
  END w_mask_in[2540]
  PIN w_mask_in[2541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.105 0.070 357.175 ;
    END
  END w_mask_in[2541]
  PIN w_mask_in[2542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.245 0.070 357.315 ;
    END
  END w_mask_in[2542]
  PIN w_mask_in[2543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.385 0.070 357.455 ;
    END
  END w_mask_in[2543]
  PIN w_mask_in[2544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.525 0.070 357.595 ;
    END
  END w_mask_in[2544]
  PIN w_mask_in[2545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.665 0.070 357.735 ;
    END
  END w_mask_in[2545]
  PIN w_mask_in[2546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.805 0.070 357.875 ;
    END
  END w_mask_in[2546]
  PIN w_mask_in[2547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 357.945 0.070 358.015 ;
    END
  END w_mask_in[2547]
  PIN w_mask_in[2548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.085 0.070 358.155 ;
    END
  END w_mask_in[2548]
  PIN w_mask_in[2549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.225 0.070 358.295 ;
    END
  END w_mask_in[2549]
  PIN w_mask_in[2550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.365 0.070 358.435 ;
    END
  END w_mask_in[2550]
  PIN w_mask_in[2551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.505 0.070 358.575 ;
    END
  END w_mask_in[2551]
  PIN w_mask_in[2552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.645 0.070 358.715 ;
    END
  END w_mask_in[2552]
  PIN w_mask_in[2553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.785 0.070 358.855 ;
    END
  END w_mask_in[2553]
  PIN w_mask_in[2554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 358.925 0.070 358.995 ;
    END
  END w_mask_in[2554]
  PIN w_mask_in[2555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.065 0.070 359.135 ;
    END
  END w_mask_in[2555]
  PIN w_mask_in[2556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.205 0.070 359.275 ;
    END
  END w_mask_in[2556]
  PIN w_mask_in[2557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.345 0.070 359.415 ;
    END
  END w_mask_in[2557]
  PIN w_mask_in[2558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.485 0.070 359.555 ;
    END
  END w_mask_in[2558]
  PIN w_mask_in[2559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.625 0.070 359.695 ;
    END
  END w_mask_in[2559]
  PIN w_mask_in[2560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.765 0.070 359.835 ;
    END
  END w_mask_in[2560]
  PIN w_mask_in[2561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.905 0.070 359.975 ;
    END
  END w_mask_in[2561]
  PIN w_mask_in[2562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.045 0.070 360.115 ;
    END
  END w_mask_in[2562]
  PIN w_mask_in[2563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.185 0.070 360.255 ;
    END
  END w_mask_in[2563]
  PIN w_mask_in[2564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.325 0.070 360.395 ;
    END
  END w_mask_in[2564]
  PIN w_mask_in[2565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.465 0.070 360.535 ;
    END
  END w_mask_in[2565]
  PIN w_mask_in[2566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.605 0.070 360.675 ;
    END
  END w_mask_in[2566]
  PIN w_mask_in[2567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.745 0.070 360.815 ;
    END
  END w_mask_in[2567]
  PIN w_mask_in[2568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 360.885 0.070 360.955 ;
    END
  END w_mask_in[2568]
  PIN w_mask_in[2569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.025 0.070 361.095 ;
    END
  END w_mask_in[2569]
  PIN w_mask_in[2570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.165 0.070 361.235 ;
    END
  END w_mask_in[2570]
  PIN w_mask_in[2571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.305 0.070 361.375 ;
    END
  END w_mask_in[2571]
  PIN w_mask_in[2572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.445 0.070 361.515 ;
    END
  END w_mask_in[2572]
  PIN w_mask_in[2573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.585 0.070 361.655 ;
    END
  END w_mask_in[2573]
  PIN w_mask_in[2574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.725 0.070 361.795 ;
    END
  END w_mask_in[2574]
  PIN w_mask_in[2575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 361.865 0.070 361.935 ;
    END
  END w_mask_in[2575]
  PIN w_mask_in[2576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.005 0.070 362.075 ;
    END
  END w_mask_in[2576]
  PIN w_mask_in[2577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.145 0.070 362.215 ;
    END
  END w_mask_in[2577]
  PIN w_mask_in[2578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.285 0.070 362.355 ;
    END
  END w_mask_in[2578]
  PIN w_mask_in[2579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.425 0.070 362.495 ;
    END
  END w_mask_in[2579]
  PIN w_mask_in[2580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.565 0.070 362.635 ;
    END
  END w_mask_in[2580]
  PIN w_mask_in[2581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.705 0.070 362.775 ;
    END
  END w_mask_in[2581]
  PIN w_mask_in[2582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.845 0.070 362.915 ;
    END
  END w_mask_in[2582]
  PIN w_mask_in[2583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.985 0.070 363.055 ;
    END
  END w_mask_in[2583]
  PIN w_mask_in[2584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.125 0.070 363.195 ;
    END
  END w_mask_in[2584]
  PIN w_mask_in[2585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.265 0.070 363.335 ;
    END
  END w_mask_in[2585]
  PIN w_mask_in[2586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.405 0.070 363.475 ;
    END
  END w_mask_in[2586]
  PIN w_mask_in[2587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.545 0.070 363.615 ;
    END
  END w_mask_in[2587]
  PIN w_mask_in[2588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.685 0.070 363.755 ;
    END
  END w_mask_in[2588]
  PIN w_mask_in[2589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.825 0.070 363.895 ;
    END
  END w_mask_in[2589]
  PIN w_mask_in[2590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 363.965 0.070 364.035 ;
    END
  END w_mask_in[2590]
  PIN w_mask_in[2591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.105 0.070 364.175 ;
    END
  END w_mask_in[2591]
  PIN w_mask_in[2592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.245 0.070 364.315 ;
    END
  END w_mask_in[2592]
  PIN w_mask_in[2593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.385 0.070 364.455 ;
    END
  END w_mask_in[2593]
  PIN w_mask_in[2594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.525 0.070 364.595 ;
    END
  END w_mask_in[2594]
  PIN w_mask_in[2595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.665 0.070 364.735 ;
    END
  END w_mask_in[2595]
  PIN w_mask_in[2596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.805 0.070 364.875 ;
    END
  END w_mask_in[2596]
  PIN w_mask_in[2597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.945 0.070 365.015 ;
    END
  END w_mask_in[2597]
  PIN w_mask_in[2598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.085 0.070 365.155 ;
    END
  END w_mask_in[2598]
  PIN w_mask_in[2599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.225 0.070 365.295 ;
    END
  END w_mask_in[2599]
  PIN w_mask_in[2600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.365 0.070 365.435 ;
    END
  END w_mask_in[2600]
  PIN w_mask_in[2601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.505 0.070 365.575 ;
    END
  END w_mask_in[2601]
  PIN w_mask_in[2602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.645 0.070 365.715 ;
    END
  END w_mask_in[2602]
  PIN w_mask_in[2603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.785 0.070 365.855 ;
    END
  END w_mask_in[2603]
  PIN w_mask_in[2604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.925 0.070 365.995 ;
    END
  END w_mask_in[2604]
  PIN w_mask_in[2605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.065 0.070 366.135 ;
    END
  END w_mask_in[2605]
  PIN w_mask_in[2606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.205 0.070 366.275 ;
    END
  END w_mask_in[2606]
  PIN w_mask_in[2607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.345 0.070 366.415 ;
    END
  END w_mask_in[2607]
  PIN w_mask_in[2608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.485 0.070 366.555 ;
    END
  END w_mask_in[2608]
  PIN w_mask_in[2609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.625 0.070 366.695 ;
    END
  END w_mask_in[2609]
  PIN w_mask_in[2610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.765 0.070 366.835 ;
    END
  END w_mask_in[2610]
  PIN w_mask_in[2611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 366.905 0.070 366.975 ;
    END
  END w_mask_in[2611]
  PIN w_mask_in[2612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.045 0.070 367.115 ;
    END
  END w_mask_in[2612]
  PIN w_mask_in[2613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.185 0.070 367.255 ;
    END
  END w_mask_in[2613]
  PIN w_mask_in[2614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.325 0.070 367.395 ;
    END
  END w_mask_in[2614]
  PIN w_mask_in[2615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.465 0.070 367.535 ;
    END
  END w_mask_in[2615]
  PIN w_mask_in[2616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.605 0.070 367.675 ;
    END
  END w_mask_in[2616]
  PIN w_mask_in[2617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.745 0.070 367.815 ;
    END
  END w_mask_in[2617]
  PIN w_mask_in[2618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.885 0.070 367.955 ;
    END
  END w_mask_in[2618]
  PIN w_mask_in[2619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.025 0.070 368.095 ;
    END
  END w_mask_in[2619]
  PIN w_mask_in[2620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.165 0.070 368.235 ;
    END
  END w_mask_in[2620]
  PIN w_mask_in[2621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.305 0.070 368.375 ;
    END
  END w_mask_in[2621]
  PIN w_mask_in[2622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.445 0.070 368.515 ;
    END
  END w_mask_in[2622]
  PIN w_mask_in[2623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.585 0.070 368.655 ;
    END
  END w_mask_in[2623]
  PIN w_mask_in[2624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.725 0.070 368.795 ;
    END
  END w_mask_in[2624]
  PIN w_mask_in[2625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 368.865 0.070 368.935 ;
    END
  END w_mask_in[2625]
  PIN w_mask_in[2626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.005 0.070 369.075 ;
    END
  END w_mask_in[2626]
  PIN w_mask_in[2627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.145 0.070 369.215 ;
    END
  END w_mask_in[2627]
  PIN w_mask_in[2628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.285 0.070 369.355 ;
    END
  END w_mask_in[2628]
  PIN w_mask_in[2629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.425 0.070 369.495 ;
    END
  END w_mask_in[2629]
  PIN w_mask_in[2630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.565 0.070 369.635 ;
    END
  END w_mask_in[2630]
  PIN w_mask_in[2631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.705 0.070 369.775 ;
    END
  END w_mask_in[2631]
  PIN w_mask_in[2632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.845 0.070 369.915 ;
    END
  END w_mask_in[2632]
  PIN w_mask_in[2633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 369.985 0.070 370.055 ;
    END
  END w_mask_in[2633]
  PIN w_mask_in[2634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.125 0.070 370.195 ;
    END
  END w_mask_in[2634]
  PIN w_mask_in[2635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.265 0.070 370.335 ;
    END
  END w_mask_in[2635]
  PIN w_mask_in[2636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.405 0.070 370.475 ;
    END
  END w_mask_in[2636]
  PIN w_mask_in[2637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.545 0.070 370.615 ;
    END
  END w_mask_in[2637]
  PIN w_mask_in[2638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.685 0.070 370.755 ;
    END
  END w_mask_in[2638]
  PIN w_mask_in[2639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.825 0.070 370.895 ;
    END
  END w_mask_in[2639]
  PIN w_mask_in[2640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.965 0.070 371.035 ;
    END
  END w_mask_in[2640]
  PIN w_mask_in[2641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.105 0.070 371.175 ;
    END
  END w_mask_in[2641]
  PIN w_mask_in[2642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.245 0.070 371.315 ;
    END
  END w_mask_in[2642]
  PIN w_mask_in[2643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.385 0.070 371.455 ;
    END
  END w_mask_in[2643]
  PIN w_mask_in[2644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.525 0.070 371.595 ;
    END
  END w_mask_in[2644]
  PIN w_mask_in[2645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.665 0.070 371.735 ;
    END
  END w_mask_in[2645]
  PIN w_mask_in[2646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.805 0.070 371.875 ;
    END
  END w_mask_in[2646]
  PIN w_mask_in[2647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 371.945 0.070 372.015 ;
    END
  END w_mask_in[2647]
  PIN w_mask_in[2648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.085 0.070 372.155 ;
    END
  END w_mask_in[2648]
  PIN w_mask_in[2649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.225 0.070 372.295 ;
    END
  END w_mask_in[2649]
  PIN w_mask_in[2650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.365 0.070 372.435 ;
    END
  END w_mask_in[2650]
  PIN w_mask_in[2651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.505 0.070 372.575 ;
    END
  END w_mask_in[2651]
  PIN w_mask_in[2652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.645 0.070 372.715 ;
    END
  END w_mask_in[2652]
  PIN w_mask_in[2653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.785 0.070 372.855 ;
    END
  END w_mask_in[2653]
  PIN w_mask_in[2654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 372.925 0.070 372.995 ;
    END
  END w_mask_in[2654]
  PIN w_mask_in[2655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.065 0.070 373.135 ;
    END
  END w_mask_in[2655]
  PIN w_mask_in[2656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.205 0.070 373.275 ;
    END
  END w_mask_in[2656]
  PIN w_mask_in[2657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.345 0.070 373.415 ;
    END
  END w_mask_in[2657]
  PIN w_mask_in[2658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.485 0.070 373.555 ;
    END
  END w_mask_in[2658]
  PIN w_mask_in[2659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.625 0.070 373.695 ;
    END
  END w_mask_in[2659]
  PIN w_mask_in[2660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.765 0.070 373.835 ;
    END
  END w_mask_in[2660]
  PIN w_mask_in[2661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.905 0.070 373.975 ;
    END
  END w_mask_in[2661]
  PIN w_mask_in[2662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.045 0.070 374.115 ;
    END
  END w_mask_in[2662]
  PIN w_mask_in[2663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.185 0.070 374.255 ;
    END
  END w_mask_in[2663]
  PIN w_mask_in[2664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.325 0.070 374.395 ;
    END
  END w_mask_in[2664]
  PIN w_mask_in[2665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.465 0.070 374.535 ;
    END
  END w_mask_in[2665]
  PIN w_mask_in[2666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.605 0.070 374.675 ;
    END
  END w_mask_in[2666]
  PIN w_mask_in[2667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.745 0.070 374.815 ;
    END
  END w_mask_in[2667]
  PIN w_mask_in[2668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 374.885 0.070 374.955 ;
    END
  END w_mask_in[2668]
  PIN w_mask_in[2669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.025 0.070 375.095 ;
    END
  END w_mask_in[2669]
  PIN w_mask_in[2670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.165 0.070 375.235 ;
    END
  END w_mask_in[2670]
  PIN w_mask_in[2671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.305 0.070 375.375 ;
    END
  END w_mask_in[2671]
  PIN w_mask_in[2672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.445 0.070 375.515 ;
    END
  END w_mask_in[2672]
  PIN w_mask_in[2673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.585 0.070 375.655 ;
    END
  END w_mask_in[2673]
  PIN w_mask_in[2674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.725 0.070 375.795 ;
    END
  END w_mask_in[2674]
  PIN w_mask_in[2675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 375.865 0.070 375.935 ;
    END
  END w_mask_in[2675]
  PIN w_mask_in[2676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.005 0.070 376.075 ;
    END
  END w_mask_in[2676]
  PIN w_mask_in[2677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.145 0.070 376.215 ;
    END
  END w_mask_in[2677]
  PIN w_mask_in[2678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.285 0.070 376.355 ;
    END
  END w_mask_in[2678]
  PIN w_mask_in[2679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.425 0.070 376.495 ;
    END
  END w_mask_in[2679]
  PIN w_mask_in[2680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.565 0.070 376.635 ;
    END
  END w_mask_in[2680]
  PIN w_mask_in[2681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.705 0.070 376.775 ;
    END
  END w_mask_in[2681]
  PIN w_mask_in[2682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.845 0.070 376.915 ;
    END
  END w_mask_in[2682]
  PIN w_mask_in[2683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.985 0.070 377.055 ;
    END
  END w_mask_in[2683]
  PIN w_mask_in[2684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.125 0.070 377.195 ;
    END
  END w_mask_in[2684]
  PIN w_mask_in[2685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.265 0.070 377.335 ;
    END
  END w_mask_in[2685]
  PIN w_mask_in[2686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.405 0.070 377.475 ;
    END
  END w_mask_in[2686]
  PIN w_mask_in[2687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.545 0.070 377.615 ;
    END
  END w_mask_in[2687]
  PIN w_mask_in[2688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.685 0.070 377.755 ;
    END
  END w_mask_in[2688]
  PIN w_mask_in[2689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.825 0.070 377.895 ;
    END
  END w_mask_in[2689]
  PIN w_mask_in[2690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 377.965 0.070 378.035 ;
    END
  END w_mask_in[2690]
  PIN w_mask_in[2691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.105 0.070 378.175 ;
    END
  END w_mask_in[2691]
  PIN w_mask_in[2692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.245 0.070 378.315 ;
    END
  END w_mask_in[2692]
  PIN w_mask_in[2693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.385 0.070 378.455 ;
    END
  END w_mask_in[2693]
  PIN w_mask_in[2694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.525 0.070 378.595 ;
    END
  END w_mask_in[2694]
  PIN w_mask_in[2695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.665 0.070 378.735 ;
    END
  END w_mask_in[2695]
  PIN w_mask_in[2696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.805 0.070 378.875 ;
    END
  END w_mask_in[2696]
  PIN w_mask_in[2697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 378.945 0.070 379.015 ;
    END
  END w_mask_in[2697]
  PIN w_mask_in[2698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.085 0.070 379.155 ;
    END
  END w_mask_in[2698]
  PIN w_mask_in[2699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.225 0.070 379.295 ;
    END
  END w_mask_in[2699]
  PIN w_mask_in[2700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.365 0.070 379.435 ;
    END
  END w_mask_in[2700]
  PIN w_mask_in[2701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.505 0.070 379.575 ;
    END
  END w_mask_in[2701]
  PIN w_mask_in[2702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.645 0.070 379.715 ;
    END
  END w_mask_in[2702]
  PIN w_mask_in[2703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.785 0.070 379.855 ;
    END
  END w_mask_in[2703]
  PIN w_mask_in[2704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 379.925 0.070 379.995 ;
    END
  END w_mask_in[2704]
  PIN w_mask_in[2705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.065 0.070 380.135 ;
    END
  END w_mask_in[2705]
  PIN w_mask_in[2706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.205 0.070 380.275 ;
    END
  END w_mask_in[2706]
  PIN w_mask_in[2707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.345 0.070 380.415 ;
    END
  END w_mask_in[2707]
  PIN w_mask_in[2708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.485 0.070 380.555 ;
    END
  END w_mask_in[2708]
  PIN w_mask_in[2709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.625 0.070 380.695 ;
    END
  END w_mask_in[2709]
  PIN w_mask_in[2710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.765 0.070 380.835 ;
    END
  END w_mask_in[2710]
  PIN w_mask_in[2711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 380.905 0.070 380.975 ;
    END
  END w_mask_in[2711]
  PIN w_mask_in[2712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.045 0.070 381.115 ;
    END
  END w_mask_in[2712]
  PIN w_mask_in[2713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.185 0.070 381.255 ;
    END
  END w_mask_in[2713]
  PIN w_mask_in[2714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.325 0.070 381.395 ;
    END
  END w_mask_in[2714]
  PIN w_mask_in[2715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.465 0.070 381.535 ;
    END
  END w_mask_in[2715]
  PIN w_mask_in[2716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.605 0.070 381.675 ;
    END
  END w_mask_in[2716]
  PIN w_mask_in[2717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.745 0.070 381.815 ;
    END
  END w_mask_in[2717]
  PIN w_mask_in[2718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.885 0.070 381.955 ;
    END
  END w_mask_in[2718]
  PIN w_mask_in[2719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.025 0.070 382.095 ;
    END
  END w_mask_in[2719]
  PIN w_mask_in[2720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.165 0.070 382.235 ;
    END
  END w_mask_in[2720]
  PIN w_mask_in[2721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.305 0.070 382.375 ;
    END
  END w_mask_in[2721]
  PIN w_mask_in[2722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.445 0.070 382.515 ;
    END
  END w_mask_in[2722]
  PIN w_mask_in[2723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.585 0.070 382.655 ;
    END
  END w_mask_in[2723]
  PIN w_mask_in[2724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.725 0.070 382.795 ;
    END
  END w_mask_in[2724]
  PIN w_mask_in[2725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 382.865 0.070 382.935 ;
    END
  END w_mask_in[2725]
  PIN w_mask_in[2726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.005 0.070 383.075 ;
    END
  END w_mask_in[2726]
  PIN w_mask_in[2727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.145 0.070 383.215 ;
    END
  END w_mask_in[2727]
  PIN w_mask_in[2728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.285 0.070 383.355 ;
    END
  END w_mask_in[2728]
  PIN w_mask_in[2729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.425 0.070 383.495 ;
    END
  END w_mask_in[2729]
  PIN w_mask_in[2730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.565 0.070 383.635 ;
    END
  END w_mask_in[2730]
  PIN w_mask_in[2731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.705 0.070 383.775 ;
    END
  END w_mask_in[2731]
  PIN w_mask_in[2732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.845 0.070 383.915 ;
    END
  END w_mask_in[2732]
  PIN w_mask_in[2733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 383.985 0.070 384.055 ;
    END
  END w_mask_in[2733]
  PIN w_mask_in[2734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.125 0.070 384.195 ;
    END
  END w_mask_in[2734]
  PIN w_mask_in[2735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.265 0.070 384.335 ;
    END
  END w_mask_in[2735]
  PIN w_mask_in[2736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.405 0.070 384.475 ;
    END
  END w_mask_in[2736]
  PIN w_mask_in[2737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.545 0.070 384.615 ;
    END
  END w_mask_in[2737]
  PIN w_mask_in[2738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.685 0.070 384.755 ;
    END
  END w_mask_in[2738]
  PIN w_mask_in[2739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.825 0.070 384.895 ;
    END
  END w_mask_in[2739]
  PIN w_mask_in[2740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.965 0.070 385.035 ;
    END
  END w_mask_in[2740]
  PIN w_mask_in[2741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.105 0.070 385.175 ;
    END
  END w_mask_in[2741]
  PIN w_mask_in[2742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.245 0.070 385.315 ;
    END
  END w_mask_in[2742]
  PIN w_mask_in[2743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.385 0.070 385.455 ;
    END
  END w_mask_in[2743]
  PIN w_mask_in[2744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.525 0.070 385.595 ;
    END
  END w_mask_in[2744]
  PIN w_mask_in[2745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.665 0.070 385.735 ;
    END
  END w_mask_in[2745]
  PIN w_mask_in[2746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.805 0.070 385.875 ;
    END
  END w_mask_in[2746]
  PIN w_mask_in[2747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 385.945 0.070 386.015 ;
    END
  END w_mask_in[2747]
  PIN w_mask_in[2748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.085 0.070 386.155 ;
    END
  END w_mask_in[2748]
  PIN w_mask_in[2749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.225 0.070 386.295 ;
    END
  END w_mask_in[2749]
  PIN w_mask_in[2750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.365 0.070 386.435 ;
    END
  END w_mask_in[2750]
  PIN w_mask_in[2751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.505 0.070 386.575 ;
    END
  END w_mask_in[2751]
  PIN w_mask_in[2752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.645 0.070 386.715 ;
    END
  END w_mask_in[2752]
  PIN w_mask_in[2753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.785 0.070 386.855 ;
    END
  END w_mask_in[2753]
  PIN w_mask_in[2754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 386.925 0.070 386.995 ;
    END
  END w_mask_in[2754]
  PIN w_mask_in[2755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.065 0.070 387.135 ;
    END
  END w_mask_in[2755]
  PIN w_mask_in[2756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.205 0.070 387.275 ;
    END
  END w_mask_in[2756]
  PIN w_mask_in[2757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.345 0.070 387.415 ;
    END
  END w_mask_in[2757]
  PIN w_mask_in[2758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.485 0.070 387.555 ;
    END
  END w_mask_in[2758]
  PIN w_mask_in[2759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.625 0.070 387.695 ;
    END
  END w_mask_in[2759]
  PIN w_mask_in[2760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.765 0.070 387.835 ;
    END
  END w_mask_in[2760]
  PIN w_mask_in[2761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.905 0.070 387.975 ;
    END
  END w_mask_in[2761]
  PIN w_mask_in[2762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.045 0.070 388.115 ;
    END
  END w_mask_in[2762]
  PIN w_mask_in[2763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.185 0.070 388.255 ;
    END
  END w_mask_in[2763]
  PIN w_mask_in[2764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.325 0.070 388.395 ;
    END
  END w_mask_in[2764]
  PIN w_mask_in[2765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.465 0.070 388.535 ;
    END
  END w_mask_in[2765]
  PIN w_mask_in[2766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.605 0.070 388.675 ;
    END
  END w_mask_in[2766]
  PIN w_mask_in[2767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.745 0.070 388.815 ;
    END
  END w_mask_in[2767]
  PIN w_mask_in[2768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 388.885 0.070 388.955 ;
    END
  END w_mask_in[2768]
  PIN w_mask_in[2769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.025 0.070 389.095 ;
    END
  END w_mask_in[2769]
  PIN w_mask_in[2770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.165 0.070 389.235 ;
    END
  END w_mask_in[2770]
  PIN w_mask_in[2771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.305 0.070 389.375 ;
    END
  END w_mask_in[2771]
  PIN w_mask_in[2772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.445 0.070 389.515 ;
    END
  END w_mask_in[2772]
  PIN w_mask_in[2773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.585 0.070 389.655 ;
    END
  END w_mask_in[2773]
  PIN w_mask_in[2774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.725 0.070 389.795 ;
    END
  END w_mask_in[2774]
  PIN w_mask_in[2775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 389.865 0.070 389.935 ;
    END
  END w_mask_in[2775]
  PIN w_mask_in[2776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.005 0.070 390.075 ;
    END
  END w_mask_in[2776]
  PIN w_mask_in[2777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.145 0.070 390.215 ;
    END
  END w_mask_in[2777]
  PIN w_mask_in[2778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.285 0.070 390.355 ;
    END
  END w_mask_in[2778]
  PIN w_mask_in[2779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.425 0.070 390.495 ;
    END
  END w_mask_in[2779]
  PIN w_mask_in[2780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.565 0.070 390.635 ;
    END
  END w_mask_in[2780]
  PIN w_mask_in[2781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.705 0.070 390.775 ;
    END
  END w_mask_in[2781]
  PIN w_mask_in[2782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.845 0.070 390.915 ;
    END
  END w_mask_in[2782]
  PIN w_mask_in[2783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.985 0.070 391.055 ;
    END
  END w_mask_in[2783]
  PIN w_mask_in[2784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.125 0.070 391.195 ;
    END
  END w_mask_in[2784]
  PIN w_mask_in[2785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.265 0.070 391.335 ;
    END
  END w_mask_in[2785]
  PIN w_mask_in[2786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.405 0.070 391.475 ;
    END
  END w_mask_in[2786]
  PIN w_mask_in[2787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.545 0.070 391.615 ;
    END
  END w_mask_in[2787]
  PIN w_mask_in[2788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.685 0.070 391.755 ;
    END
  END w_mask_in[2788]
  PIN w_mask_in[2789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.825 0.070 391.895 ;
    END
  END w_mask_in[2789]
  PIN w_mask_in[2790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 391.965 0.070 392.035 ;
    END
  END w_mask_in[2790]
  PIN w_mask_in[2791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.105 0.070 392.175 ;
    END
  END w_mask_in[2791]
  PIN w_mask_in[2792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.245 0.070 392.315 ;
    END
  END w_mask_in[2792]
  PIN w_mask_in[2793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.385 0.070 392.455 ;
    END
  END w_mask_in[2793]
  PIN w_mask_in[2794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.525 0.070 392.595 ;
    END
  END w_mask_in[2794]
  PIN w_mask_in[2795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.665 0.070 392.735 ;
    END
  END w_mask_in[2795]
  PIN w_mask_in[2796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.805 0.070 392.875 ;
    END
  END w_mask_in[2796]
  PIN w_mask_in[2797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 392.945 0.070 393.015 ;
    END
  END w_mask_in[2797]
  PIN w_mask_in[2798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.085 0.070 393.155 ;
    END
  END w_mask_in[2798]
  PIN w_mask_in[2799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.225 0.070 393.295 ;
    END
  END w_mask_in[2799]
  PIN w_mask_in[2800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.365 0.070 393.435 ;
    END
  END w_mask_in[2800]
  PIN w_mask_in[2801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.505 0.070 393.575 ;
    END
  END w_mask_in[2801]
  PIN w_mask_in[2802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.645 0.070 393.715 ;
    END
  END w_mask_in[2802]
  PIN w_mask_in[2803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.785 0.070 393.855 ;
    END
  END w_mask_in[2803]
  PIN w_mask_in[2804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.925 0.070 393.995 ;
    END
  END w_mask_in[2804]
  PIN w_mask_in[2805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.065 0.070 394.135 ;
    END
  END w_mask_in[2805]
  PIN w_mask_in[2806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.205 0.070 394.275 ;
    END
  END w_mask_in[2806]
  PIN w_mask_in[2807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.345 0.070 394.415 ;
    END
  END w_mask_in[2807]
  PIN w_mask_in[2808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.485 0.070 394.555 ;
    END
  END w_mask_in[2808]
  PIN w_mask_in[2809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.625 0.070 394.695 ;
    END
  END w_mask_in[2809]
  PIN w_mask_in[2810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.765 0.070 394.835 ;
    END
  END w_mask_in[2810]
  PIN w_mask_in[2811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 394.905 0.070 394.975 ;
    END
  END w_mask_in[2811]
  PIN w_mask_in[2812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.045 0.070 395.115 ;
    END
  END w_mask_in[2812]
  PIN w_mask_in[2813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.185 0.070 395.255 ;
    END
  END w_mask_in[2813]
  PIN w_mask_in[2814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.325 0.070 395.395 ;
    END
  END w_mask_in[2814]
  PIN w_mask_in[2815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.465 0.070 395.535 ;
    END
  END w_mask_in[2815]
  PIN w_mask_in[2816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.605 0.070 395.675 ;
    END
  END w_mask_in[2816]
  PIN w_mask_in[2817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.745 0.070 395.815 ;
    END
  END w_mask_in[2817]
  PIN w_mask_in[2818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 395.885 0.070 395.955 ;
    END
  END w_mask_in[2818]
  PIN w_mask_in[2819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.025 0.070 396.095 ;
    END
  END w_mask_in[2819]
  PIN w_mask_in[2820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.165 0.070 396.235 ;
    END
  END w_mask_in[2820]
  PIN w_mask_in[2821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.305 0.070 396.375 ;
    END
  END w_mask_in[2821]
  PIN w_mask_in[2822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.445 0.070 396.515 ;
    END
  END w_mask_in[2822]
  PIN w_mask_in[2823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.585 0.070 396.655 ;
    END
  END w_mask_in[2823]
  PIN w_mask_in[2824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.725 0.070 396.795 ;
    END
  END w_mask_in[2824]
  PIN w_mask_in[2825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.865 0.070 396.935 ;
    END
  END w_mask_in[2825]
  PIN w_mask_in[2826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.005 0.070 397.075 ;
    END
  END w_mask_in[2826]
  PIN w_mask_in[2827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.145 0.070 397.215 ;
    END
  END w_mask_in[2827]
  PIN w_mask_in[2828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.285 0.070 397.355 ;
    END
  END w_mask_in[2828]
  PIN w_mask_in[2829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.425 0.070 397.495 ;
    END
  END w_mask_in[2829]
  PIN w_mask_in[2830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.565 0.070 397.635 ;
    END
  END w_mask_in[2830]
  PIN w_mask_in[2831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.705 0.070 397.775 ;
    END
  END w_mask_in[2831]
  PIN w_mask_in[2832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.845 0.070 397.915 ;
    END
  END w_mask_in[2832]
  PIN w_mask_in[2833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 397.985 0.070 398.055 ;
    END
  END w_mask_in[2833]
  PIN w_mask_in[2834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.125 0.070 398.195 ;
    END
  END w_mask_in[2834]
  PIN w_mask_in[2835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.265 0.070 398.335 ;
    END
  END w_mask_in[2835]
  PIN w_mask_in[2836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.405 0.070 398.475 ;
    END
  END w_mask_in[2836]
  PIN w_mask_in[2837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.545 0.070 398.615 ;
    END
  END w_mask_in[2837]
  PIN w_mask_in[2838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.685 0.070 398.755 ;
    END
  END w_mask_in[2838]
  PIN w_mask_in[2839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.825 0.070 398.895 ;
    END
  END w_mask_in[2839]
  PIN w_mask_in[2840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 398.965 0.070 399.035 ;
    END
  END w_mask_in[2840]
  PIN w_mask_in[2841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.105 0.070 399.175 ;
    END
  END w_mask_in[2841]
  PIN w_mask_in[2842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.245 0.070 399.315 ;
    END
  END w_mask_in[2842]
  PIN w_mask_in[2843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.385 0.070 399.455 ;
    END
  END w_mask_in[2843]
  PIN w_mask_in[2844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.525 0.070 399.595 ;
    END
  END w_mask_in[2844]
  PIN w_mask_in[2845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.665 0.070 399.735 ;
    END
  END w_mask_in[2845]
  PIN w_mask_in[2846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.805 0.070 399.875 ;
    END
  END w_mask_in[2846]
  PIN w_mask_in[2847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.945 0.070 400.015 ;
    END
  END w_mask_in[2847]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.525 0.070 504.595 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.665 0.070 504.735 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.805 0.070 504.875 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 504.945 0.070 505.015 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.085 0.070 505.155 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.225 0.070 505.295 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.365 0.070 505.435 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.505 0.070 505.575 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.645 0.070 505.715 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.785 0.070 505.855 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.925 0.070 505.995 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.065 0.070 506.135 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.205 0.070 506.275 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.345 0.070 506.415 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.485 0.070 506.555 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.625 0.070 506.695 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.765 0.070 506.835 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 506.905 0.070 506.975 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.045 0.070 507.115 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.185 0.070 507.255 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.325 0.070 507.395 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.465 0.070 507.535 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.605 0.070 507.675 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.745 0.070 507.815 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 507.885 0.070 507.955 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.025 0.070 508.095 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.165 0.070 508.235 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.305 0.070 508.375 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.445 0.070 508.515 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.585 0.070 508.655 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.725 0.070 508.795 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.865 0.070 508.935 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.005 0.070 509.075 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.145 0.070 509.215 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.285 0.070 509.355 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.425 0.070 509.495 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.565 0.070 509.635 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.705 0.070 509.775 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.845 0.070 509.915 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 509.985 0.070 510.055 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.125 0.070 510.195 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.265 0.070 510.335 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.405 0.070 510.475 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.545 0.070 510.615 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.685 0.070 510.755 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.825 0.070 510.895 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.965 0.070 511.035 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.105 0.070 511.175 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.245 0.070 511.315 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.385 0.070 511.455 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.525 0.070 511.595 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.665 0.070 511.735 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.805 0.070 511.875 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 511.945 0.070 512.015 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.085 0.070 512.155 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.225 0.070 512.295 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.365 0.070 512.435 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.505 0.070 512.575 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.645 0.070 512.715 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.785 0.070 512.855 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 512.925 0.070 512.995 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.065 0.070 513.135 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.205 0.070 513.275 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.345 0.070 513.415 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.485 0.070 513.555 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.625 0.070 513.695 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.765 0.070 513.835 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.905 0.070 513.975 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.045 0.070 514.115 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.185 0.070 514.255 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.325 0.070 514.395 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.465 0.070 514.535 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.605 0.070 514.675 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.745 0.070 514.815 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 514.885 0.070 514.955 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.025 0.070 515.095 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.165 0.070 515.235 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.305 0.070 515.375 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.445 0.070 515.515 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.585 0.070 515.655 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.725 0.070 515.795 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 515.865 0.070 515.935 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.005 0.070 516.075 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.145 0.070 516.215 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.285 0.070 516.355 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.425 0.070 516.495 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.565 0.070 516.635 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.705 0.070 516.775 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.845 0.070 516.915 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.985 0.070 517.055 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.125 0.070 517.195 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.265 0.070 517.335 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.405 0.070 517.475 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.545 0.070 517.615 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.685 0.070 517.755 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.825 0.070 517.895 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 517.965 0.070 518.035 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.105 0.070 518.175 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.245 0.070 518.315 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.385 0.070 518.455 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.525 0.070 518.595 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.665 0.070 518.735 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.805 0.070 518.875 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 518.945 0.070 519.015 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.085 0.070 519.155 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.225 0.070 519.295 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.365 0.070 519.435 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.505 0.070 519.575 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.645 0.070 519.715 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.785 0.070 519.855 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.925 0.070 519.995 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.065 0.070 520.135 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.205 0.070 520.275 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.345 0.070 520.415 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.485 0.070 520.555 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.625 0.070 520.695 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.765 0.070 520.835 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 520.905 0.070 520.975 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.045 0.070 521.115 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.185 0.070 521.255 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.325 0.070 521.395 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.465 0.070 521.535 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.605 0.070 521.675 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.745 0.070 521.815 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 521.885 0.070 521.955 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.025 0.070 522.095 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.165 0.070 522.235 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.305 0.070 522.375 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.445 0.070 522.515 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.585 0.070 522.655 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.725 0.070 522.795 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.865 0.070 522.935 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.005 0.070 523.075 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.145 0.070 523.215 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.285 0.070 523.355 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.425 0.070 523.495 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.565 0.070 523.635 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.705 0.070 523.775 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.845 0.070 523.915 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 523.985 0.070 524.055 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.125 0.070 524.195 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.265 0.070 524.335 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.405 0.070 524.475 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.545 0.070 524.615 ;
    END
  END rd_out[143]
  PIN rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.685 0.070 524.755 ;
    END
  END rd_out[144]
  PIN rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.825 0.070 524.895 ;
    END
  END rd_out[145]
  PIN rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 524.965 0.070 525.035 ;
    END
  END rd_out[146]
  PIN rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.105 0.070 525.175 ;
    END
  END rd_out[147]
  PIN rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.245 0.070 525.315 ;
    END
  END rd_out[148]
  PIN rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.385 0.070 525.455 ;
    END
  END rd_out[149]
  PIN rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.525 0.070 525.595 ;
    END
  END rd_out[150]
  PIN rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.665 0.070 525.735 ;
    END
  END rd_out[151]
  PIN rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.805 0.070 525.875 ;
    END
  END rd_out[152]
  PIN rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.945 0.070 526.015 ;
    END
  END rd_out[153]
  PIN rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.085 0.070 526.155 ;
    END
  END rd_out[154]
  PIN rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.225 0.070 526.295 ;
    END
  END rd_out[155]
  PIN rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.365 0.070 526.435 ;
    END
  END rd_out[156]
  PIN rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.505 0.070 526.575 ;
    END
  END rd_out[157]
  PIN rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.645 0.070 526.715 ;
    END
  END rd_out[158]
  PIN rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.785 0.070 526.855 ;
    END
  END rd_out[159]
  PIN rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 526.925 0.070 526.995 ;
    END
  END rd_out[160]
  PIN rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.065 0.070 527.135 ;
    END
  END rd_out[161]
  PIN rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.205 0.070 527.275 ;
    END
  END rd_out[162]
  PIN rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.345 0.070 527.415 ;
    END
  END rd_out[163]
  PIN rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.485 0.070 527.555 ;
    END
  END rd_out[164]
  PIN rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.625 0.070 527.695 ;
    END
  END rd_out[165]
  PIN rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.765 0.070 527.835 ;
    END
  END rd_out[166]
  PIN rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 527.905 0.070 527.975 ;
    END
  END rd_out[167]
  PIN rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.045 0.070 528.115 ;
    END
  END rd_out[168]
  PIN rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.185 0.070 528.255 ;
    END
  END rd_out[169]
  PIN rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.325 0.070 528.395 ;
    END
  END rd_out[170]
  PIN rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.465 0.070 528.535 ;
    END
  END rd_out[171]
  PIN rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.605 0.070 528.675 ;
    END
  END rd_out[172]
  PIN rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.745 0.070 528.815 ;
    END
  END rd_out[173]
  PIN rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.885 0.070 528.955 ;
    END
  END rd_out[174]
  PIN rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.025 0.070 529.095 ;
    END
  END rd_out[175]
  PIN rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.165 0.070 529.235 ;
    END
  END rd_out[176]
  PIN rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.305 0.070 529.375 ;
    END
  END rd_out[177]
  PIN rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.445 0.070 529.515 ;
    END
  END rd_out[178]
  PIN rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.585 0.070 529.655 ;
    END
  END rd_out[179]
  PIN rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.725 0.070 529.795 ;
    END
  END rd_out[180]
  PIN rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 529.865 0.070 529.935 ;
    END
  END rd_out[181]
  PIN rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.005 0.070 530.075 ;
    END
  END rd_out[182]
  PIN rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.145 0.070 530.215 ;
    END
  END rd_out[183]
  PIN rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.285 0.070 530.355 ;
    END
  END rd_out[184]
  PIN rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.425 0.070 530.495 ;
    END
  END rd_out[185]
  PIN rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.565 0.070 530.635 ;
    END
  END rd_out[186]
  PIN rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.705 0.070 530.775 ;
    END
  END rd_out[187]
  PIN rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.845 0.070 530.915 ;
    END
  END rd_out[188]
  PIN rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 530.985 0.070 531.055 ;
    END
  END rd_out[189]
  PIN rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.125 0.070 531.195 ;
    END
  END rd_out[190]
  PIN rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.265 0.070 531.335 ;
    END
  END rd_out[191]
  PIN rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.405 0.070 531.475 ;
    END
  END rd_out[192]
  PIN rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.545 0.070 531.615 ;
    END
  END rd_out[193]
  PIN rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.685 0.070 531.755 ;
    END
  END rd_out[194]
  PIN rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.825 0.070 531.895 ;
    END
  END rd_out[195]
  PIN rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.965 0.070 532.035 ;
    END
  END rd_out[196]
  PIN rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.105 0.070 532.175 ;
    END
  END rd_out[197]
  PIN rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.245 0.070 532.315 ;
    END
  END rd_out[198]
  PIN rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.385 0.070 532.455 ;
    END
  END rd_out[199]
  PIN rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.525 0.070 532.595 ;
    END
  END rd_out[200]
  PIN rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.665 0.070 532.735 ;
    END
  END rd_out[201]
  PIN rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.805 0.070 532.875 ;
    END
  END rd_out[202]
  PIN rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 532.945 0.070 533.015 ;
    END
  END rd_out[203]
  PIN rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.085 0.070 533.155 ;
    END
  END rd_out[204]
  PIN rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.225 0.070 533.295 ;
    END
  END rd_out[205]
  PIN rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.365 0.070 533.435 ;
    END
  END rd_out[206]
  PIN rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.505 0.070 533.575 ;
    END
  END rd_out[207]
  PIN rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.645 0.070 533.715 ;
    END
  END rd_out[208]
  PIN rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.785 0.070 533.855 ;
    END
  END rd_out[209]
  PIN rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 533.925 0.070 533.995 ;
    END
  END rd_out[210]
  PIN rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.065 0.070 534.135 ;
    END
  END rd_out[211]
  PIN rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.205 0.070 534.275 ;
    END
  END rd_out[212]
  PIN rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.345 0.070 534.415 ;
    END
  END rd_out[213]
  PIN rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.485 0.070 534.555 ;
    END
  END rd_out[214]
  PIN rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.625 0.070 534.695 ;
    END
  END rd_out[215]
  PIN rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.765 0.070 534.835 ;
    END
  END rd_out[216]
  PIN rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.905 0.070 534.975 ;
    END
  END rd_out[217]
  PIN rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.045 0.070 535.115 ;
    END
  END rd_out[218]
  PIN rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.185 0.070 535.255 ;
    END
  END rd_out[219]
  PIN rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.325 0.070 535.395 ;
    END
  END rd_out[220]
  PIN rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.465 0.070 535.535 ;
    END
  END rd_out[221]
  PIN rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.605 0.070 535.675 ;
    END
  END rd_out[222]
  PIN rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.745 0.070 535.815 ;
    END
  END rd_out[223]
  PIN rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 535.885 0.070 535.955 ;
    END
  END rd_out[224]
  PIN rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.025 0.070 536.095 ;
    END
  END rd_out[225]
  PIN rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.165 0.070 536.235 ;
    END
  END rd_out[226]
  PIN rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.305 0.070 536.375 ;
    END
  END rd_out[227]
  PIN rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.445 0.070 536.515 ;
    END
  END rd_out[228]
  PIN rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.585 0.070 536.655 ;
    END
  END rd_out[229]
  PIN rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.725 0.070 536.795 ;
    END
  END rd_out[230]
  PIN rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 536.865 0.070 536.935 ;
    END
  END rd_out[231]
  PIN rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.005 0.070 537.075 ;
    END
  END rd_out[232]
  PIN rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.145 0.070 537.215 ;
    END
  END rd_out[233]
  PIN rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.285 0.070 537.355 ;
    END
  END rd_out[234]
  PIN rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.425 0.070 537.495 ;
    END
  END rd_out[235]
  PIN rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.565 0.070 537.635 ;
    END
  END rd_out[236]
  PIN rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.705 0.070 537.775 ;
    END
  END rd_out[237]
  PIN rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.845 0.070 537.915 ;
    END
  END rd_out[238]
  PIN rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.985 0.070 538.055 ;
    END
  END rd_out[239]
  PIN rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.125 0.070 538.195 ;
    END
  END rd_out[240]
  PIN rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.265 0.070 538.335 ;
    END
  END rd_out[241]
  PIN rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.405 0.070 538.475 ;
    END
  END rd_out[242]
  PIN rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.545 0.070 538.615 ;
    END
  END rd_out[243]
  PIN rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.685 0.070 538.755 ;
    END
  END rd_out[244]
  PIN rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.825 0.070 538.895 ;
    END
  END rd_out[245]
  PIN rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 538.965 0.070 539.035 ;
    END
  END rd_out[246]
  PIN rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.105 0.070 539.175 ;
    END
  END rd_out[247]
  PIN rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.245 0.070 539.315 ;
    END
  END rd_out[248]
  PIN rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.385 0.070 539.455 ;
    END
  END rd_out[249]
  PIN rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.525 0.070 539.595 ;
    END
  END rd_out[250]
  PIN rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.665 0.070 539.735 ;
    END
  END rd_out[251]
  PIN rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.805 0.070 539.875 ;
    END
  END rd_out[252]
  PIN rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 539.945 0.070 540.015 ;
    END
  END rd_out[253]
  PIN rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.085 0.070 540.155 ;
    END
  END rd_out[254]
  PIN rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.225 0.070 540.295 ;
    END
  END rd_out[255]
  PIN rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.365 0.070 540.435 ;
    END
  END rd_out[256]
  PIN rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.505 0.070 540.575 ;
    END
  END rd_out[257]
  PIN rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.645 0.070 540.715 ;
    END
  END rd_out[258]
  PIN rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.785 0.070 540.855 ;
    END
  END rd_out[259]
  PIN rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.925 0.070 540.995 ;
    END
  END rd_out[260]
  PIN rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.065 0.070 541.135 ;
    END
  END rd_out[261]
  PIN rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.205 0.070 541.275 ;
    END
  END rd_out[262]
  PIN rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.345 0.070 541.415 ;
    END
  END rd_out[263]
  PIN rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.485 0.070 541.555 ;
    END
  END rd_out[264]
  PIN rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.625 0.070 541.695 ;
    END
  END rd_out[265]
  PIN rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.765 0.070 541.835 ;
    END
  END rd_out[266]
  PIN rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 541.905 0.070 541.975 ;
    END
  END rd_out[267]
  PIN rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.045 0.070 542.115 ;
    END
  END rd_out[268]
  PIN rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.185 0.070 542.255 ;
    END
  END rd_out[269]
  PIN rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.325 0.070 542.395 ;
    END
  END rd_out[270]
  PIN rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.465 0.070 542.535 ;
    END
  END rd_out[271]
  PIN rd_out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.605 0.070 542.675 ;
    END
  END rd_out[272]
  PIN rd_out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.745 0.070 542.815 ;
    END
  END rd_out[273]
  PIN rd_out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 542.885 0.070 542.955 ;
    END
  END rd_out[274]
  PIN rd_out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.025 0.070 543.095 ;
    END
  END rd_out[275]
  PIN rd_out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.165 0.070 543.235 ;
    END
  END rd_out[276]
  PIN rd_out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.305 0.070 543.375 ;
    END
  END rd_out[277]
  PIN rd_out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.445 0.070 543.515 ;
    END
  END rd_out[278]
  PIN rd_out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.585 0.070 543.655 ;
    END
  END rd_out[279]
  PIN rd_out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.725 0.070 543.795 ;
    END
  END rd_out[280]
  PIN rd_out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.865 0.070 543.935 ;
    END
  END rd_out[281]
  PIN rd_out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.005 0.070 544.075 ;
    END
  END rd_out[282]
  PIN rd_out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.145 0.070 544.215 ;
    END
  END rd_out[283]
  PIN rd_out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.285 0.070 544.355 ;
    END
  END rd_out[284]
  PIN rd_out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.425 0.070 544.495 ;
    END
  END rd_out[285]
  PIN rd_out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.565 0.070 544.635 ;
    END
  END rd_out[286]
  PIN rd_out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.705 0.070 544.775 ;
    END
  END rd_out[287]
  PIN rd_out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.845 0.070 544.915 ;
    END
  END rd_out[288]
  PIN rd_out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 544.985 0.070 545.055 ;
    END
  END rd_out[289]
  PIN rd_out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.125 0.070 545.195 ;
    END
  END rd_out[290]
  PIN rd_out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.265 0.070 545.335 ;
    END
  END rd_out[291]
  PIN rd_out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.405 0.070 545.475 ;
    END
  END rd_out[292]
  PIN rd_out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.545 0.070 545.615 ;
    END
  END rd_out[293]
  PIN rd_out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.685 0.070 545.755 ;
    END
  END rd_out[294]
  PIN rd_out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.825 0.070 545.895 ;
    END
  END rd_out[295]
  PIN rd_out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 545.965 0.070 546.035 ;
    END
  END rd_out[296]
  PIN rd_out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.105 0.070 546.175 ;
    END
  END rd_out[297]
  PIN rd_out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.245 0.070 546.315 ;
    END
  END rd_out[298]
  PIN rd_out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.385 0.070 546.455 ;
    END
  END rd_out[299]
  PIN rd_out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.525 0.070 546.595 ;
    END
  END rd_out[300]
  PIN rd_out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.665 0.070 546.735 ;
    END
  END rd_out[301]
  PIN rd_out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.805 0.070 546.875 ;
    END
  END rd_out[302]
  PIN rd_out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.945 0.070 547.015 ;
    END
  END rd_out[303]
  PIN rd_out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.085 0.070 547.155 ;
    END
  END rd_out[304]
  PIN rd_out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.225 0.070 547.295 ;
    END
  END rd_out[305]
  PIN rd_out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.365 0.070 547.435 ;
    END
  END rd_out[306]
  PIN rd_out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.505 0.070 547.575 ;
    END
  END rd_out[307]
  PIN rd_out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.645 0.070 547.715 ;
    END
  END rd_out[308]
  PIN rd_out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.785 0.070 547.855 ;
    END
  END rd_out[309]
  PIN rd_out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 547.925 0.070 547.995 ;
    END
  END rd_out[310]
  PIN rd_out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.065 0.070 548.135 ;
    END
  END rd_out[311]
  PIN rd_out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.205 0.070 548.275 ;
    END
  END rd_out[312]
  PIN rd_out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.345 0.070 548.415 ;
    END
  END rd_out[313]
  PIN rd_out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.485 0.070 548.555 ;
    END
  END rd_out[314]
  PIN rd_out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.625 0.070 548.695 ;
    END
  END rd_out[315]
  PIN rd_out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.765 0.070 548.835 ;
    END
  END rd_out[316]
  PIN rd_out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 548.905 0.070 548.975 ;
    END
  END rd_out[317]
  PIN rd_out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.045 0.070 549.115 ;
    END
  END rd_out[318]
  PIN rd_out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.185 0.070 549.255 ;
    END
  END rd_out[319]
  PIN rd_out[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.325 0.070 549.395 ;
    END
  END rd_out[320]
  PIN rd_out[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.465 0.070 549.535 ;
    END
  END rd_out[321]
  PIN rd_out[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.605 0.070 549.675 ;
    END
  END rd_out[322]
  PIN rd_out[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.745 0.070 549.815 ;
    END
  END rd_out[323]
  PIN rd_out[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.885 0.070 549.955 ;
    END
  END rd_out[324]
  PIN rd_out[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.025 0.070 550.095 ;
    END
  END rd_out[325]
  PIN rd_out[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.165 0.070 550.235 ;
    END
  END rd_out[326]
  PIN rd_out[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.305 0.070 550.375 ;
    END
  END rd_out[327]
  PIN rd_out[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.445 0.070 550.515 ;
    END
  END rd_out[328]
  PIN rd_out[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.585 0.070 550.655 ;
    END
  END rd_out[329]
  PIN rd_out[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.725 0.070 550.795 ;
    END
  END rd_out[330]
  PIN rd_out[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 550.865 0.070 550.935 ;
    END
  END rd_out[331]
  PIN rd_out[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.005 0.070 551.075 ;
    END
  END rd_out[332]
  PIN rd_out[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.145 0.070 551.215 ;
    END
  END rd_out[333]
  PIN rd_out[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.285 0.070 551.355 ;
    END
  END rd_out[334]
  PIN rd_out[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.425 0.070 551.495 ;
    END
  END rd_out[335]
  PIN rd_out[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.565 0.070 551.635 ;
    END
  END rd_out[336]
  PIN rd_out[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.705 0.070 551.775 ;
    END
  END rd_out[337]
  PIN rd_out[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.845 0.070 551.915 ;
    END
  END rd_out[338]
  PIN rd_out[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 551.985 0.070 552.055 ;
    END
  END rd_out[339]
  PIN rd_out[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.125 0.070 552.195 ;
    END
  END rd_out[340]
  PIN rd_out[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.265 0.070 552.335 ;
    END
  END rd_out[341]
  PIN rd_out[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.405 0.070 552.475 ;
    END
  END rd_out[342]
  PIN rd_out[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.545 0.070 552.615 ;
    END
  END rd_out[343]
  PIN rd_out[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.685 0.070 552.755 ;
    END
  END rd_out[344]
  PIN rd_out[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.825 0.070 552.895 ;
    END
  END rd_out[345]
  PIN rd_out[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.965 0.070 553.035 ;
    END
  END rd_out[346]
  PIN rd_out[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.105 0.070 553.175 ;
    END
  END rd_out[347]
  PIN rd_out[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.245 0.070 553.315 ;
    END
  END rd_out[348]
  PIN rd_out[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.385 0.070 553.455 ;
    END
  END rd_out[349]
  PIN rd_out[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.525 0.070 553.595 ;
    END
  END rd_out[350]
  PIN rd_out[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.665 0.070 553.735 ;
    END
  END rd_out[351]
  PIN rd_out[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.805 0.070 553.875 ;
    END
  END rd_out[352]
  PIN rd_out[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 553.945 0.070 554.015 ;
    END
  END rd_out[353]
  PIN rd_out[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.085 0.070 554.155 ;
    END
  END rd_out[354]
  PIN rd_out[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.225 0.070 554.295 ;
    END
  END rd_out[355]
  PIN rd_out[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.365 0.070 554.435 ;
    END
  END rd_out[356]
  PIN rd_out[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.505 0.070 554.575 ;
    END
  END rd_out[357]
  PIN rd_out[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.645 0.070 554.715 ;
    END
  END rd_out[358]
  PIN rd_out[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.785 0.070 554.855 ;
    END
  END rd_out[359]
  PIN rd_out[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 554.925 0.070 554.995 ;
    END
  END rd_out[360]
  PIN rd_out[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.065 0.070 555.135 ;
    END
  END rd_out[361]
  PIN rd_out[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.205 0.070 555.275 ;
    END
  END rd_out[362]
  PIN rd_out[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.345 0.070 555.415 ;
    END
  END rd_out[363]
  PIN rd_out[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.485 0.070 555.555 ;
    END
  END rd_out[364]
  PIN rd_out[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.625 0.070 555.695 ;
    END
  END rd_out[365]
  PIN rd_out[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.765 0.070 555.835 ;
    END
  END rd_out[366]
  PIN rd_out[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.905 0.070 555.975 ;
    END
  END rd_out[367]
  PIN rd_out[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.045 0.070 556.115 ;
    END
  END rd_out[368]
  PIN rd_out[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.185 0.070 556.255 ;
    END
  END rd_out[369]
  PIN rd_out[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.325 0.070 556.395 ;
    END
  END rd_out[370]
  PIN rd_out[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.465 0.070 556.535 ;
    END
  END rd_out[371]
  PIN rd_out[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.605 0.070 556.675 ;
    END
  END rd_out[372]
  PIN rd_out[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.745 0.070 556.815 ;
    END
  END rd_out[373]
  PIN rd_out[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 556.885 0.070 556.955 ;
    END
  END rd_out[374]
  PIN rd_out[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.025 0.070 557.095 ;
    END
  END rd_out[375]
  PIN rd_out[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.165 0.070 557.235 ;
    END
  END rd_out[376]
  PIN rd_out[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.305 0.070 557.375 ;
    END
  END rd_out[377]
  PIN rd_out[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.445 0.070 557.515 ;
    END
  END rd_out[378]
  PIN rd_out[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.585 0.070 557.655 ;
    END
  END rd_out[379]
  PIN rd_out[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.725 0.070 557.795 ;
    END
  END rd_out[380]
  PIN rd_out[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 557.865 0.070 557.935 ;
    END
  END rd_out[381]
  PIN rd_out[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.005 0.070 558.075 ;
    END
  END rd_out[382]
  PIN rd_out[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.145 0.070 558.215 ;
    END
  END rd_out[383]
  PIN rd_out[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.285 0.070 558.355 ;
    END
  END rd_out[384]
  PIN rd_out[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.425 0.070 558.495 ;
    END
  END rd_out[385]
  PIN rd_out[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.565 0.070 558.635 ;
    END
  END rd_out[386]
  PIN rd_out[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.705 0.070 558.775 ;
    END
  END rd_out[387]
  PIN rd_out[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.845 0.070 558.915 ;
    END
  END rd_out[388]
  PIN rd_out[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.985 0.070 559.055 ;
    END
  END rd_out[389]
  PIN rd_out[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.125 0.070 559.195 ;
    END
  END rd_out[390]
  PIN rd_out[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.265 0.070 559.335 ;
    END
  END rd_out[391]
  PIN rd_out[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.405 0.070 559.475 ;
    END
  END rd_out[392]
  PIN rd_out[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.545 0.070 559.615 ;
    END
  END rd_out[393]
  PIN rd_out[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.685 0.070 559.755 ;
    END
  END rd_out[394]
  PIN rd_out[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.825 0.070 559.895 ;
    END
  END rd_out[395]
  PIN rd_out[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 559.965 0.070 560.035 ;
    END
  END rd_out[396]
  PIN rd_out[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.105 0.070 560.175 ;
    END
  END rd_out[397]
  PIN rd_out[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.245 0.070 560.315 ;
    END
  END rd_out[398]
  PIN rd_out[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.385 0.070 560.455 ;
    END
  END rd_out[399]
  PIN rd_out[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.525 0.070 560.595 ;
    END
  END rd_out[400]
  PIN rd_out[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.665 0.070 560.735 ;
    END
  END rd_out[401]
  PIN rd_out[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.805 0.070 560.875 ;
    END
  END rd_out[402]
  PIN rd_out[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.945 0.070 561.015 ;
    END
  END rd_out[403]
  PIN rd_out[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.085 0.070 561.155 ;
    END
  END rd_out[404]
  PIN rd_out[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.225 0.070 561.295 ;
    END
  END rd_out[405]
  PIN rd_out[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.365 0.070 561.435 ;
    END
  END rd_out[406]
  PIN rd_out[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.505 0.070 561.575 ;
    END
  END rd_out[407]
  PIN rd_out[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.645 0.070 561.715 ;
    END
  END rd_out[408]
  PIN rd_out[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.785 0.070 561.855 ;
    END
  END rd_out[409]
  PIN rd_out[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 561.925 0.070 561.995 ;
    END
  END rd_out[410]
  PIN rd_out[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.065 0.070 562.135 ;
    END
  END rd_out[411]
  PIN rd_out[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.205 0.070 562.275 ;
    END
  END rd_out[412]
  PIN rd_out[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.345 0.070 562.415 ;
    END
  END rd_out[413]
  PIN rd_out[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.485 0.070 562.555 ;
    END
  END rd_out[414]
  PIN rd_out[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.625 0.070 562.695 ;
    END
  END rd_out[415]
  PIN rd_out[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.765 0.070 562.835 ;
    END
  END rd_out[416]
  PIN rd_out[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 562.905 0.070 562.975 ;
    END
  END rd_out[417]
  PIN rd_out[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.045 0.070 563.115 ;
    END
  END rd_out[418]
  PIN rd_out[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.185 0.070 563.255 ;
    END
  END rd_out[419]
  PIN rd_out[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.325 0.070 563.395 ;
    END
  END rd_out[420]
  PIN rd_out[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.465 0.070 563.535 ;
    END
  END rd_out[421]
  PIN rd_out[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.605 0.070 563.675 ;
    END
  END rd_out[422]
  PIN rd_out[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.745 0.070 563.815 ;
    END
  END rd_out[423]
  PIN rd_out[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.885 0.070 563.955 ;
    END
  END rd_out[424]
  PIN rd_out[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.025 0.070 564.095 ;
    END
  END rd_out[425]
  PIN rd_out[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.165 0.070 564.235 ;
    END
  END rd_out[426]
  PIN rd_out[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.305 0.070 564.375 ;
    END
  END rd_out[427]
  PIN rd_out[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.445 0.070 564.515 ;
    END
  END rd_out[428]
  PIN rd_out[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.585 0.070 564.655 ;
    END
  END rd_out[429]
  PIN rd_out[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.725 0.070 564.795 ;
    END
  END rd_out[430]
  PIN rd_out[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 564.865 0.070 564.935 ;
    END
  END rd_out[431]
  PIN rd_out[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.005 0.070 565.075 ;
    END
  END rd_out[432]
  PIN rd_out[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.145 0.070 565.215 ;
    END
  END rd_out[433]
  PIN rd_out[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.285 0.070 565.355 ;
    END
  END rd_out[434]
  PIN rd_out[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.425 0.070 565.495 ;
    END
  END rd_out[435]
  PIN rd_out[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.565 0.070 565.635 ;
    END
  END rd_out[436]
  PIN rd_out[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.705 0.070 565.775 ;
    END
  END rd_out[437]
  PIN rd_out[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.845 0.070 565.915 ;
    END
  END rd_out[438]
  PIN rd_out[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 565.985 0.070 566.055 ;
    END
  END rd_out[439]
  PIN rd_out[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.125 0.070 566.195 ;
    END
  END rd_out[440]
  PIN rd_out[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.265 0.070 566.335 ;
    END
  END rd_out[441]
  PIN rd_out[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.405 0.070 566.475 ;
    END
  END rd_out[442]
  PIN rd_out[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.545 0.070 566.615 ;
    END
  END rd_out[443]
  PIN rd_out[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.685 0.070 566.755 ;
    END
  END rd_out[444]
  PIN rd_out[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.825 0.070 566.895 ;
    END
  END rd_out[445]
  PIN rd_out[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.965 0.070 567.035 ;
    END
  END rd_out[446]
  PIN rd_out[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.105 0.070 567.175 ;
    END
  END rd_out[447]
  PIN rd_out[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.245 0.070 567.315 ;
    END
  END rd_out[448]
  PIN rd_out[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.385 0.070 567.455 ;
    END
  END rd_out[449]
  PIN rd_out[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.525 0.070 567.595 ;
    END
  END rd_out[450]
  PIN rd_out[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.665 0.070 567.735 ;
    END
  END rd_out[451]
  PIN rd_out[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.805 0.070 567.875 ;
    END
  END rd_out[452]
  PIN rd_out[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 567.945 0.070 568.015 ;
    END
  END rd_out[453]
  PIN rd_out[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.085 0.070 568.155 ;
    END
  END rd_out[454]
  PIN rd_out[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.225 0.070 568.295 ;
    END
  END rd_out[455]
  PIN rd_out[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.365 0.070 568.435 ;
    END
  END rd_out[456]
  PIN rd_out[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.505 0.070 568.575 ;
    END
  END rd_out[457]
  PIN rd_out[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.645 0.070 568.715 ;
    END
  END rd_out[458]
  PIN rd_out[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.785 0.070 568.855 ;
    END
  END rd_out[459]
  PIN rd_out[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 568.925 0.070 568.995 ;
    END
  END rd_out[460]
  PIN rd_out[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.065 0.070 569.135 ;
    END
  END rd_out[461]
  PIN rd_out[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.205 0.070 569.275 ;
    END
  END rd_out[462]
  PIN rd_out[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.345 0.070 569.415 ;
    END
  END rd_out[463]
  PIN rd_out[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.485 0.070 569.555 ;
    END
  END rd_out[464]
  PIN rd_out[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.625 0.070 569.695 ;
    END
  END rd_out[465]
  PIN rd_out[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.765 0.070 569.835 ;
    END
  END rd_out[466]
  PIN rd_out[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 569.905 0.070 569.975 ;
    END
  END rd_out[467]
  PIN rd_out[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.045 0.070 570.115 ;
    END
  END rd_out[468]
  PIN rd_out[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.185 0.070 570.255 ;
    END
  END rd_out[469]
  PIN rd_out[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.325 0.070 570.395 ;
    END
  END rd_out[470]
  PIN rd_out[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.465 0.070 570.535 ;
    END
  END rd_out[471]
  PIN rd_out[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.605 0.070 570.675 ;
    END
  END rd_out[472]
  PIN rd_out[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.745 0.070 570.815 ;
    END
  END rd_out[473]
  PIN rd_out[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 570.885 0.070 570.955 ;
    END
  END rd_out[474]
  PIN rd_out[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.025 0.070 571.095 ;
    END
  END rd_out[475]
  PIN rd_out[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.165 0.070 571.235 ;
    END
  END rd_out[476]
  PIN rd_out[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.305 0.070 571.375 ;
    END
  END rd_out[477]
  PIN rd_out[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.445 0.070 571.515 ;
    END
  END rd_out[478]
  PIN rd_out[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.585 0.070 571.655 ;
    END
  END rd_out[479]
  PIN rd_out[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.725 0.070 571.795 ;
    END
  END rd_out[480]
  PIN rd_out[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.865 0.070 571.935 ;
    END
  END rd_out[481]
  PIN rd_out[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.005 0.070 572.075 ;
    END
  END rd_out[482]
  PIN rd_out[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.145 0.070 572.215 ;
    END
  END rd_out[483]
  PIN rd_out[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.285 0.070 572.355 ;
    END
  END rd_out[484]
  PIN rd_out[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.425 0.070 572.495 ;
    END
  END rd_out[485]
  PIN rd_out[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.565 0.070 572.635 ;
    END
  END rd_out[486]
  PIN rd_out[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.705 0.070 572.775 ;
    END
  END rd_out[487]
  PIN rd_out[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.845 0.070 572.915 ;
    END
  END rd_out[488]
  PIN rd_out[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 572.985 0.070 573.055 ;
    END
  END rd_out[489]
  PIN rd_out[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.125 0.070 573.195 ;
    END
  END rd_out[490]
  PIN rd_out[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.265 0.070 573.335 ;
    END
  END rd_out[491]
  PIN rd_out[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.405 0.070 573.475 ;
    END
  END rd_out[492]
  PIN rd_out[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.545 0.070 573.615 ;
    END
  END rd_out[493]
  PIN rd_out[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.685 0.070 573.755 ;
    END
  END rd_out[494]
  PIN rd_out[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.825 0.070 573.895 ;
    END
  END rd_out[495]
  PIN rd_out[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 573.965 0.070 574.035 ;
    END
  END rd_out[496]
  PIN rd_out[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.105 0.070 574.175 ;
    END
  END rd_out[497]
  PIN rd_out[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.245 0.070 574.315 ;
    END
  END rd_out[498]
  PIN rd_out[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.385 0.070 574.455 ;
    END
  END rd_out[499]
  PIN rd_out[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.525 0.070 574.595 ;
    END
  END rd_out[500]
  PIN rd_out[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.665 0.070 574.735 ;
    END
  END rd_out[501]
  PIN rd_out[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.805 0.070 574.875 ;
    END
  END rd_out[502]
  PIN rd_out[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.945 0.070 575.015 ;
    END
  END rd_out[503]
  PIN rd_out[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.085 0.070 575.155 ;
    END
  END rd_out[504]
  PIN rd_out[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.225 0.070 575.295 ;
    END
  END rd_out[505]
  PIN rd_out[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.365 0.070 575.435 ;
    END
  END rd_out[506]
  PIN rd_out[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.505 0.070 575.575 ;
    END
  END rd_out[507]
  PIN rd_out[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.645 0.070 575.715 ;
    END
  END rd_out[508]
  PIN rd_out[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.785 0.070 575.855 ;
    END
  END rd_out[509]
  PIN rd_out[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 575.925 0.070 575.995 ;
    END
  END rd_out[510]
  PIN rd_out[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.065 0.070 576.135 ;
    END
  END rd_out[511]
  PIN rd_out[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.205 0.070 576.275 ;
    END
  END rd_out[512]
  PIN rd_out[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.345 0.070 576.415 ;
    END
  END rd_out[513]
  PIN rd_out[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.485 0.070 576.555 ;
    END
  END rd_out[514]
  PIN rd_out[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.625 0.070 576.695 ;
    END
  END rd_out[515]
  PIN rd_out[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.765 0.070 576.835 ;
    END
  END rd_out[516]
  PIN rd_out[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 576.905 0.070 576.975 ;
    END
  END rd_out[517]
  PIN rd_out[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.045 0.070 577.115 ;
    END
  END rd_out[518]
  PIN rd_out[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.185 0.070 577.255 ;
    END
  END rd_out[519]
  PIN rd_out[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.325 0.070 577.395 ;
    END
  END rd_out[520]
  PIN rd_out[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.465 0.070 577.535 ;
    END
  END rd_out[521]
  PIN rd_out[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.605 0.070 577.675 ;
    END
  END rd_out[522]
  PIN rd_out[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.745 0.070 577.815 ;
    END
  END rd_out[523]
  PIN rd_out[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.885 0.070 577.955 ;
    END
  END rd_out[524]
  PIN rd_out[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.025 0.070 578.095 ;
    END
  END rd_out[525]
  PIN rd_out[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.165 0.070 578.235 ;
    END
  END rd_out[526]
  PIN rd_out[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.305 0.070 578.375 ;
    END
  END rd_out[527]
  PIN rd_out[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.445 0.070 578.515 ;
    END
  END rd_out[528]
  PIN rd_out[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.585 0.070 578.655 ;
    END
  END rd_out[529]
  PIN rd_out[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.725 0.070 578.795 ;
    END
  END rd_out[530]
  PIN rd_out[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 578.865 0.070 578.935 ;
    END
  END rd_out[531]
  PIN rd_out[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.005 0.070 579.075 ;
    END
  END rd_out[532]
  PIN rd_out[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.145 0.070 579.215 ;
    END
  END rd_out[533]
  PIN rd_out[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.285 0.070 579.355 ;
    END
  END rd_out[534]
  PIN rd_out[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.425 0.070 579.495 ;
    END
  END rd_out[535]
  PIN rd_out[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.565 0.070 579.635 ;
    END
  END rd_out[536]
  PIN rd_out[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.705 0.070 579.775 ;
    END
  END rd_out[537]
  PIN rd_out[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.845 0.070 579.915 ;
    END
  END rd_out[538]
  PIN rd_out[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 579.985 0.070 580.055 ;
    END
  END rd_out[539]
  PIN rd_out[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.125 0.070 580.195 ;
    END
  END rd_out[540]
  PIN rd_out[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.265 0.070 580.335 ;
    END
  END rd_out[541]
  PIN rd_out[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.405 0.070 580.475 ;
    END
  END rd_out[542]
  PIN rd_out[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.545 0.070 580.615 ;
    END
  END rd_out[543]
  PIN rd_out[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.685 0.070 580.755 ;
    END
  END rd_out[544]
  PIN rd_out[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.825 0.070 580.895 ;
    END
  END rd_out[545]
  PIN rd_out[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.965 0.070 581.035 ;
    END
  END rd_out[546]
  PIN rd_out[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.105 0.070 581.175 ;
    END
  END rd_out[547]
  PIN rd_out[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.245 0.070 581.315 ;
    END
  END rd_out[548]
  PIN rd_out[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.385 0.070 581.455 ;
    END
  END rd_out[549]
  PIN rd_out[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.525 0.070 581.595 ;
    END
  END rd_out[550]
  PIN rd_out[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.665 0.070 581.735 ;
    END
  END rd_out[551]
  PIN rd_out[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.805 0.070 581.875 ;
    END
  END rd_out[552]
  PIN rd_out[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 581.945 0.070 582.015 ;
    END
  END rd_out[553]
  PIN rd_out[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.085 0.070 582.155 ;
    END
  END rd_out[554]
  PIN rd_out[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.225 0.070 582.295 ;
    END
  END rd_out[555]
  PIN rd_out[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.365 0.070 582.435 ;
    END
  END rd_out[556]
  PIN rd_out[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.505 0.070 582.575 ;
    END
  END rd_out[557]
  PIN rd_out[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.645 0.070 582.715 ;
    END
  END rd_out[558]
  PIN rd_out[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.785 0.070 582.855 ;
    END
  END rd_out[559]
  PIN rd_out[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 582.925 0.070 582.995 ;
    END
  END rd_out[560]
  PIN rd_out[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.065 0.070 583.135 ;
    END
  END rd_out[561]
  PIN rd_out[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.205 0.070 583.275 ;
    END
  END rd_out[562]
  PIN rd_out[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.345 0.070 583.415 ;
    END
  END rd_out[563]
  PIN rd_out[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.485 0.070 583.555 ;
    END
  END rd_out[564]
  PIN rd_out[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.625 0.070 583.695 ;
    END
  END rd_out[565]
  PIN rd_out[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.765 0.070 583.835 ;
    END
  END rd_out[566]
  PIN rd_out[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.905 0.070 583.975 ;
    END
  END rd_out[567]
  PIN rd_out[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.045 0.070 584.115 ;
    END
  END rd_out[568]
  PIN rd_out[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.185 0.070 584.255 ;
    END
  END rd_out[569]
  PIN rd_out[570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.325 0.070 584.395 ;
    END
  END rd_out[570]
  PIN rd_out[571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.465 0.070 584.535 ;
    END
  END rd_out[571]
  PIN rd_out[572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.605 0.070 584.675 ;
    END
  END rd_out[572]
  PIN rd_out[573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.745 0.070 584.815 ;
    END
  END rd_out[573]
  PIN rd_out[574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 584.885 0.070 584.955 ;
    END
  END rd_out[574]
  PIN rd_out[575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.025 0.070 585.095 ;
    END
  END rd_out[575]
  PIN rd_out[576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.165 0.070 585.235 ;
    END
  END rd_out[576]
  PIN rd_out[577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.305 0.070 585.375 ;
    END
  END rd_out[577]
  PIN rd_out[578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.445 0.070 585.515 ;
    END
  END rd_out[578]
  PIN rd_out[579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.585 0.070 585.655 ;
    END
  END rd_out[579]
  PIN rd_out[580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.725 0.070 585.795 ;
    END
  END rd_out[580]
  PIN rd_out[581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 585.865 0.070 585.935 ;
    END
  END rd_out[581]
  PIN rd_out[582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.005 0.070 586.075 ;
    END
  END rd_out[582]
  PIN rd_out[583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.145 0.070 586.215 ;
    END
  END rd_out[583]
  PIN rd_out[584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.285 0.070 586.355 ;
    END
  END rd_out[584]
  PIN rd_out[585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.425 0.070 586.495 ;
    END
  END rd_out[585]
  PIN rd_out[586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.565 0.070 586.635 ;
    END
  END rd_out[586]
  PIN rd_out[587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.705 0.070 586.775 ;
    END
  END rd_out[587]
  PIN rd_out[588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.845 0.070 586.915 ;
    END
  END rd_out[588]
  PIN rd_out[589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.985 0.070 587.055 ;
    END
  END rd_out[589]
  PIN rd_out[590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.125 0.070 587.195 ;
    END
  END rd_out[590]
  PIN rd_out[591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.265 0.070 587.335 ;
    END
  END rd_out[591]
  PIN rd_out[592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.405 0.070 587.475 ;
    END
  END rd_out[592]
  PIN rd_out[593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.545 0.070 587.615 ;
    END
  END rd_out[593]
  PIN rd_out[594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.685 0.070 587.755 ;
    END
  END rd_out[594]
  PIN rd_out[595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.825 0.070 587.895 ;
    END
  END rd_out[595]
  PIN rd_out[596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 587.965 0.070 588.035 ;
    END
  END rd_out[596]
  PIN rd_out[597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.105 0.070 588.175 ;
    END
  END rd_out[597]
  PIN rd_out[598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.245 0.070 588.315 ;
    END
  END rd_out[598]
  PIN rd_out[599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.385 0.070 588.455 ;
    END
  END rd_out[599]
  PIN rd_out[600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.525 0.070 588.595 ;
    END
  END rd_out[600]
  PIN rd_out[601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.665 0.070 588.735 ;
    END
  END rd_out[601]
  PIN rd_out[602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.805 0.070 588.875 ;
    END
  END rd_out[602]
  PIN rd_out[603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 588.945 0.070 589.015 ;
    END
  END rd_out[603]
  PIN rd_out[604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.085 0.070 589.155 ;
    END
  END rd_out[604]
  PIN rd_out[605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.225 0.070 589.295 ;
    END
  END rd_out[605]
  PIN rd_out[606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.365 0.070 589.435 ;
    END
  END rd_out[606]
  PIN rd_out[607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.505 0.070 589.575 ;
    END
  END rd_out[607]
  PIN rd_out[608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.645 0.070 589.715 ;
    END
  END rd_out[608]
  PIN rd_out[609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.785 0.070 589.855 ;
    END
  END rd_out[609]
  PIN rd_out[610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.925 0.070 589.995 ;
    END
  END rd_out[610]
  PIN rd_out[611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.065 0.070 590.135 ;
    END
  END rd_out[611]
  PIN rd_out[612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.205 0.070 590.275 ;
    END
  END rd_out[612]
  PIN rd_out[613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.345 0.070 590.415 ;
    END
  END rd_out[613]
  PIN rd_out[614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.485 0.070 590.555 ;
    END
  END rd_out[614]
  PIN rd_out[615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.625 0.070 590.695 ;
    END
  END rd_out[615]
  PIN rd_out[616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.765 0.070 590.835 ;
    END
  END rd_out[616]
  PIN rd_out[617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 590.905 0.070 590.975 ;
    END
  END rd_out[617]
  PIN rd_out[618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.045 0.070 591.115 ;
    END
  END rd_out[618]
  PIN rd_out[619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.185 0.070 591.255 ;
    END
  END rd_out[619]
  PIN rd_out[620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.325 0.070 591.395 ;
    END
  END rd_out[620]
  PIN rd_out[621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.465 0.070 591.535 ;
    END
  END rd_out[621]
  PIN rd_out[622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.605 0.070 591.675 ;
    END
  END rd_out[622]
  PIN rd_out[623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.745 0.070 591.815 ;
    END
  END rd_out[623]
  PIN rd_out[624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 591.885 0.070 591.955 ;
    END
  END rd_out[624]
  PIN rd_out[625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.025 0.070 592.095 ;
    END
  END rd_out[625]
  PIN rd_out[626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.165 0.070 592.235 ;
    END
  END rd_out[626]
  PIN rd_out[627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.305 0.070 592.375 ;
    END
  END rd_out[627]
  PIN rd_out[628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.445 0.070 592.515 ;
    END
  END rd_out[628]
  PIN rd_out[629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.585 0.070 592.655 ;
    END
  END rd_out[629]
  PIN rd_out[630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.725 0.070 592.795 ;
    END
  END rd_out[630]
  PIN rd_out[631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.865 0.070 592.935 ;
    END
  END rd_out[631]
  PIN rd_out[632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.005 0.070 593.075 ;
    END
  END rd_out[632]
  PIN rd_out[633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.145 0.070 593.215 ;
    END
  END rd_out[633]
  PIN rd_out[634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.285 0.070 593.355 ;
    END
  END rd_out[634]
  PIN rd_out[635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.425 0.070 593.495 ;
    END
  END rd_out[635]
  PIN rd_out[636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.565 0.070 593.635 ;
    END
  END rd_out[636]
  PIN rd_out[637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.705 0.070 593.775 ;
    END
  END rd_out[637]
  PIN rd_out[638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.845 0.070 593.915 ;
    END
  END rd_out[638]
  PIN rd_out[639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 593.985 0.070 594.055 ;
    END
  END rd_out[639]
  PIN rd_out[640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.125 0.070 594.195 ;
    END
  END rd_out[640]
  PIN rd_out[641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.265 0.070 594.335 ;
    END
  END rd_out[641]
  PIN rd_out[642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.405 0.070 594.475 ;
    END
  END rd_out[642]
  PIN rd_out[643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.545 0.070 594.615 ;
    END
  END rd_out[643]
  PIN rd_out[644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.685 0.070 594.755 ;
    END
  END rd_out[644]
  PIN rd_out[645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.825 0.070 594.895 ;
    END
  END rd_out[645]
  PIN rd_out[646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 594.965 0.070 595.035 ;
    END
  END rd_out[646]
  PIN rd_out[647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.105 0.070 595.175 ;
    END
  END rd_out[647]
  PIN rd_out[648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.245 0.070 595.315 ;
    END
  END rd_out[648]
  PIN rd_out[649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.385 0.070 595.455 ;
    END
  END rd_out[649]
  PIN rd_out[650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.525 0.070 595.595 ;
    END
  END rd_out[650]
  PIN rd_out[651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.665 0.070 595.735 ;
    END
  END rd_out[651]
  PIN rd_out[652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.805 0.070 595.875 ;
    END
  END rd_out[652]
  PIN rd_out[653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.945 0.070 596.015 ;
    END
  END rd_out[653]
  PIN rd_out[654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.085 0.070 596.155 ;
    END
  END rd_out[654]
  PIN rd_out[655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.225 0.070 596.295 ;
    END
  END rd_out[655]
  PIN rd_out[656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.365 0.070 596.435 ;
    END
  END rd_out[656]
  PIN rd_out[657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.505 0.070 596.575 ;
    END
  END rd_out[657]
  PIN rd_out[658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.645 0.070 596.715 ;
    END
  END rd_out[658]
  PIN rd_out[659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.785 0.070 596.855 ;
    END
  END rd_out[659]
  PIN rd_out[660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 596.925 0.070 596.995 ;
    END
  END rd_out[660]
  PIN rd_out[661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.065 0.070 597.135 ;
    END
  END rd_out[661]
  PIN rd_out[662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.205 0.070 597.275 ;
    END
  END rd_out[662]
  PIN rd_out[663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.345 0.070 597.415 ;
    END
  END rd_out[663]
  PIN rd_out[664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.485 0.070 597.555 ;
    END
  END rd_out[664]
  PIN rd_out[665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.625 0.070 597.695 ;
    END
  END rd_out[665]
  PIN rd_out[666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.765 0.070 597.835 ;
    END
  END rd_out[666]
  PIN rd_out[667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 597.905 0.070 597.975 ;
    END
  END rd_out[667]
  PIN rd_out[668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.045 0.070 598.115 ;
    END
  END rd_out[668]
  PIN rd_out[669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.185 0.070 598.255 ;
    END
  END rd_out[669]
  PIN rd_out[670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.325 0.070 598.395 ;
    END
  END rd_out[670]
  PIN rd_out[671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.465 0.070 598.535 ;
    END
  END rd_out[671]
  PIN rd_out[672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.605 0.070 598.675 ;
    END
  END rd_out[672]
  PIN rd_out[673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.745 0.070 598.815 ;
    END
  END rd_out[673]
  PIN rd_out[674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.885 0.070 598.955 ;
    END
  END rd_out[674]
  PIN rd_out[675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.025 0.070 599.095 ;
    END
  END rd_out[675]
  PIN rd_out[676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.165 0.070 599.235 ;
    END
  END rd_out[676]
  PIN rd_out[677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.305 0.070 599.375 ;
    END
  END rd_out[677]
  PIN rd_out[678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.445 0.070 599.515 ;
    END
  END rd_out[678]
  PIN rd_out[679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.585 0.070 599.655 ;
    END
  END rd_out[679]
  PIN rd_out[680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.725 0.070 599.795 ;
    END
  END rd_out[680]
  PIN rd_out[681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 599.865 0.070 599.935 ;
    END
  END rd_out[681]
  PIN rd_out[682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.005 0.070 600.075 ;
    END
  END rd_out[682]
  PIN rd_out[683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.145 0.070 600.215 ;
    END
  END rd_out[683]
  PIN rd_out[684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.285 0.070 600.355 ;
    END
  END rd_out[684]
  PIN rd_out[685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.425 0.070 600.495 ;
    END
  END rd_out[685]
  PIN rd_out[686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.565 0.070 600.635 ;
    END
  END rd_out[686]
  PIN rd_out[687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.705 0.070 600.775 ;
    END
  END rd_out[687]
  PIN rd_out[688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.845 0.070 600.915 ;
    END
  END rd_out[688]
  PIN rd_out[689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 600.985 0.070 601.055 ;
    END
  END rd_out[689]
  PIN rd_out[690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.125 0.070 601.195 ;
    END
  END rd_out[690]
  PIN rd_out[691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.265 0.070 601.335 ;
    END
  END rd_out[691]
  PIN rd_out[692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.405 0.070 601.475 ;
    END
  END rd_out[692]
  PIN rd_out[693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.545 0.070 601.615 ;
    END
  END rd_out[693]
  PIN rd_out[694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.685 0.070 601.755 ;
    END
  END rd_out[694]
  PIN rd_out[695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.825 0.070 601.895 ;
    END
  END rd_out[695]
  PIN rd_out[696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.965 0.070 602.035 ;
    END
  END rd_out[696]
  PIN rd_out[697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.105 0.070 602.175 ;
    END
  END rd_out[697]
  PIN rd_out[698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.245 0.070 602.315 ;
    END
  END rd_out[698]
  PIN rd_out[699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.385 0.070 602.455 ;
    END
  END rd_out[699]
  PIN rd_out[700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.525 0.070 602.595 ;
    END
  END rd_out[700]
  PIN rd_out[701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.665 0.070 602.735 ;
    END
  END rd_out[701]
  PIN rd_out[702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.805 0.070 602.875 ;
    END
  END rd_out[702]
  PIN rd_out[703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 602.945 0.070 603.015 ;
    END
  END rd_out[703]
  PIN rd_out[704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.085 0.070 603.155 ;
    END
  END rd_out[704]
  PIN rd_out[705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.225 0.070 603.295 ;
    END
  END rd_out[705]
  PIN rd_out[706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.365 0.070 603.435 ;
    END
  END rd_out[706]
  PIN rd_out[707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.505 0.070 603.575 ;
    END
  END rd_out[707]
  PIN rd_out[708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.645 0.070 603.715 ;
    END
  END rd_out[708]
  PIN rd_out[709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.785 0.070 603.855 ;
    END
  END rd_out[709]
  PIN rd_out[710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 603.925 0.070 603.995 ;
    END
  END rd_out[710]
  PIN rd_out[711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.065 0.070 604.135 ;
    END
  END rd_out[711]
  PIN rd_out[712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.205 0.070 604.275 ;
    END
  END rd_out[712]
  PIN rd_out[713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.345 0.070 604.415 ;
    END
  END rd_out[713]
  PIN rd_out[714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.485 0.070 604.555 ;
    END
  END rd_out[714]
  PIN rd_out[715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.625 0.070 604.695 ;
    END
  END rd_out[715]
  PIN rd_out[716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.765 0.070 604.835 ;
    END
  END rd_out[716]
  PIN rd_out[717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.905 0.070 604.975 ;
    END
  END rd_out[717]
  PIN rd_out[718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.045 0.070 605.115 ;
    END
  END rd_out[718]
  PIN rd_out[719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.185 0.070 605.255 ;
    END
  END rd_out[719]
  PIN rd_out[720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.325 0.070 605.395 ;
    END
  END rd_out[720]
  PIN rd_out[721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.465 0.070 605.535 ;
    END
  END rd_out[721]
  PIN rd_out[722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.605 0.070 605.675 ;
    END
  END rd_out[722]
  PIN rd_out[723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.745 0.070 605.815 ;
    END
  END rd_out[723]
  PIN rd_out[724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 605.885 0.070 605.955 ;
    END
  END rd_out[724]
  PIN rd_out[725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.025 0.070 606.095 ;
    END
  END rd_out[725]
  PIN rd_out[726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.165 0.070 606.235 ;
    END
  END rd_out[726]
  PIN rd_out[727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.305 0.070 606.375 ;
    END
  END rd_out[727]
  PIN rd_out[728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.445 0.070 606.515 ;
    END
  END rd_out[728]
  PIN rd_out[729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.585 0.070 606.655 ;
    END
  END rd_out[729]
  PIN rd_out[730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.725 0.070 606.795 ;
    END
  END rd_out[730]
  PIN rd_out[731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 606.865 0.070 606.935 ;
    END
  END rd_out[731]
  PIN rd_out[732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.005 0.070 607.075 ;
    END
  END rd_out[732]
  PIN rd_out[733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.145 0.070 607.215 ;
    END
  END rd_out[733]
  PIN rd_out[734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.285 0.070 607.355 ;
    END
  END rd_out[734]
  PIN rd_out[735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.425 0.070 607.495 ;
    END
  END rd_out[735]
  PIN rd_out[736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.565 0.070 607.635 ;
    END
  END rd_out[736]
  PIN rd_out[737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.705 0.070 607.775 ;
    END
  END rd_out[737]
  PIN rd_out[738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.845 0.070 607.915 ;
    END
  END rd_out[738]
  PIN rd_out[739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.985 0.070 608.055 ;
    END
  END rd_out[739]
  PIN rd_out[740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.125 0.070 608.195 ;
    END
  END rd_out[740]
  PIN rd_out[741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.265 0.070 608.335 ;
    END
  END rd_out[741]
  PIN rd_out[742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.405 0.070 608.475 ;
    END
  END rd_out[742]
  PIN rd_out[743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.545 0.070 608.615 ;
    END
  END rd_out[743]
  PIN rd_out[744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.685 0.070 608.755 ;
    END
  END rd_out[744]
  PIN rd_out[745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.825 0.070 608.895 ;
    END
  END rd_out[745]
  PIN rd_out[746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 608.965 0.070 609.035 ;
    END
  END rd_out[746]
  PIN rd_out[747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.105 0.070 609.175 ;
    END
  END rd_out[747]
  PIN rd_out[748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.245 0.070 609.315 ;
    END
  END rd_out[748]
  PIN rd_out[749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.385 0.070 609.455 ;
    END
  END rd_out[749]
  PIN rd_out[750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.525 0.070 609.595 ;
    END
  END rd_out[750]
  PIN rd_out[751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.665 0.070 609.735 ;
    END
  END rd_out[751]
  PIN rd_out[752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.805 0.070 609.875 ;
    END
  END rd_out[752]
  PIN rd_out[753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.945 0.070 610.015 ;
    END
  END rd_out[753]
  PIN rd_out[754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.085 0.070 610.155 ;
    END
  END rd_out[754]
  PIN rd_out[755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.225 0.070 610.295 ;
    END
  END rd_out[755]
  PIN rd_out[756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.365 0.070 610.435 ;
    END
  END rd_out[756]
  PIN rd_out[757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.505 0.070 610.575 ;
    END
  END rd_out[757]
  PIN rd_out[758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.645 0.070 610.715 ;
    END
  END rd_out[758]
  PIN rd_out[759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.785 0.070 610.855 ;
    END
  END rd_out[759]
  PIN rd_out[760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 610.925 0.070 610.995 ;
    END
  END rd_out[760]
  PIN rd_out[761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.065 0.070 611.135 ;
    END
  END rd_out[761]
  PIN rd_out[762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.205 0.070 611.275 ;
    END
  END rd_out[762]
  PIN rd_out[763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.345 0.070 611.415 ;
    END
  END rd_out[763]
  PIN rd_out[764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.485 0.070 611.555 ;
    END
  END rd_out[764]
  PIN rd_out[765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.625 0.070 611.695 ;
    END
  END rd_out[765]
  PIN rd_out[766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.765 0.070 611.835 ;
    END
  END rd_out[766]
  PIN rd_out[767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 611.905 0.070 611.975 ;
    END
  END rd_out[767]
  PIN rd_out[768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.045 0.070 612.115 ;
    END
  END rd_out[768]
  PIN rd_out[769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.185 0.070 612.255 ;
    END
  END rd_out[769]
  PIN rd_out[770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.325 0.070 612.395 ;
    END
  END rd_out[770]
  PIN rd_out[771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.465 0.070 612.535 ;
    END
  END rd_out[771]
  PIN rd_out[772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.605 0.070 612.675 ;
    END
  END rd_out[772]
  PIN rd_out[773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.745 0.070 612.815 ;
    END
  END rd_out[773]
  PIN rd_out[774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 612.885 0.070 612.955 ;
    END
  END rd_out[774]
  PIN rd_out[775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.025 0.070 613.095 ;
    END
  END rd_out[775]
  PIN rd_out[776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.165 0.070 613.235 ;
    END
  END rd_out[776]
  PIN rd_out[777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.305 0.070 613.375 ;
    END
  END rd_out[777]
  PIN rd_out[778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.445 0.070 613.515 ;
    END
  END rd_out[778]
  PIN rd_out[779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.585 0.070 613.655 ;
    END
  END rd_out[779]
  PIN rd_out[780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.725 0.070 613.795 ;
    END
  END rd_out[780]
  PIN rd_out[781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 613.865 0.070 613.935 ;
    END
  END rd_out[781]
  PIN rd_out[782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.005 0.070 614.075 ;
    END
  END rd_out[782]
  PIN rd_out[783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.145 0.070 614.215 ;
    END
  END rd_out[783]
  PIN rd_out[784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.285 0.070 614.355 ;
    END
  END rd_out[784]
  PIN rd_out[785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.425 0.070 614.495 ;
    END
  END rd_out[785]
  PIN rd_out[786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.565 0.070 614.635 ;
    END
  END rd_out[786]
  PIN rd_out[787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.705 0.070 614.775 ;
    END
  END rd_out[787]
  PIN rd_out[788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.845 0.070 614.915 ;
    END
  END rd_out[788]
  PIN rd_out[789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.985 0.070 615.055 ;
    END
  END rd_out[789]
  PIN rd_out[790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.125 0.070 615.195 ;
    END
  END rd_out[790]
  PIN rd_out[791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.265 0.070 615.335 ;
    END
  END rd_out[791]
  PIN rd_out[792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.405 0.070 615.475 ;
    END
  END rd_out[792]
  PIN rd_out[793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.545 0.070 615.615 ;
    END
  END rd_out[793]
  PIN rd_out[794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.685 0.070 615.755 ;
    END
  END rd_out[794]
  PIN rd_out[795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.825 0.070 615.895 ;
    END
  END rd_out[795]
  PIN rd_out[796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 615.965 0.070 616.035 ;
    END
  END rd_out[796]
  PIN rd_out[797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.105 0.070 616.175 ;
    END
  END rd_out[797]
  PIN rd_out[798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.245 0.070 616.315 ;
    END
  END rd_out[798]
  PIN rd_out[799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.385 0.070 616.455 ;
    END
  END rd_out[799]
  PIN rd_out[800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.525 0.070 616.595 ;
    END
  END rd_out[800]
  PIN rd_out[801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.665 0.070 616.735 ;
    END
  END rd_out[801]
  PIN rd_out[802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.805 0.070 616.875 ;
    END
  END rd_out[802]
  PIN rd_out[803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 616.945 0.070 617.015 ;
    END
  END rd_out[803]
  PIN rd_out[804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.085 0.070 617.155 ;
    END
  END rd_out[804]
  PIN rd_out[805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.225 0.070 617.295 ;
    END
  END rd_out[805]
  PIN rd_out[806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.365 0.070 617.435 ;
    END
  END rd_out[806]
  PIN rd_out[807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.505 0.070 617.575 ;
    END
  END rd_out[807]
  PIN rd_out[808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.645 0.070 617.715 ;
    END
  END rd_out[808]
  PIN rd_out[809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.785 0.070 617.855 ;
    END
  END rd_out[809]
  PIN rd_out[810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.925 0.070 617.995 ;
    END
  END rd_out[810]
  PIN rd_out[811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.065 0.070 618.135 ;
    END
  END rd_out[811]
  PIN rd_out[812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.205 0.070 618.275 ;
    END
  END rd_out[812]
  PIN rd_out[813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.345 0.070 618.415 ;
    END
  END rd_out[813]
  PIN rd_out[814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.485 0.070 618.555 ;
    END
  END rd_out[814]
  PIN rd_out[815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.625 0.070 618.695 ;
    END
  END rd_out[815]
  PIN rd_out[816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.765 0.070 618.835 ;
    END
  END rd_out[816]
  PIN rd_out[817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 618.905 0.070 618.975 ;
    END
  END rd_out[817]
  PIN rd_out[818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.045 0.070 619.115 ;
    END
  END rd_out[818]
  PIN rd_out[819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.185 0.070 619.255 ;
    END
  END rd_out[819]
  PIN rd_out[820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.325 0.070 619.395 ;
    END
  END rd_out[820]
  PIN rd_out[821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.465 0.070 619.535 ;
    END
  END rd_out[821]
  PIN rd_out[822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.605 0.070 619.675 ;
    END
  END rd_out[822]
  PIN rd_out[823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.745 0.070 619.815 ;
    END
  END rd_out[823]
  PIN rd_out[824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 619.885 0.070 619.955 ;
    END
  END rd_out[824]
  PIN rd_out[825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.025 0.070 620.095 ;
    END
  END rd_out[825]
  PIN rd_out[826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.165 0.070 620.235 ;
    END
  END rd_out[826]
  PIN rd_out[827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.305 0.070 620.375 ;
    END
  END rd_out[827]
  PIN rd_out[828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.445 0.070 620.515 ;
    END
  END rd_out[828]
  PIN rd_out[829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.585 0.070 620.655 ;
    END
  END rd_out[829]
  PIN rd_out[830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.725 0.070 620.795 ;
    END
  END rd_out[830]
  PIN rd_out[831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.865 0.070 620.935 ;
    END
  END rd_out[831]
  PIN rd_out[832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.005 0.070 621.075 ;
    END
  END rd_out[832]
  PIN rd_out[833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.145 0.070 621.215 ;
    END
  END rd_out[833]
  PIN rd_out[834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.285 0.070 621.355 ;
    END
  END rd_out[834]
  PIN rd_out[835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.425 0.070 621.495 ;
    END
  END rd_out[835]
  PIN rd_out[836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.565 0.070 621.635 ;
    END
  END rd_out[836]
  PIN rd_out[837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.705 0.070 621.775 ;
    END
  END rd_out[837]
  PIN rd_out[838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.845 0.070 621.915 ;
    END
  END rd_out[838]
  PIN rd_out[839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 621.985 0.070 622.055 ;
    END
  END rd_out[839]
  PIN rd_out[840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.125 0.070 622.195 ;
    END
  END rd_out[840]
  PIN rd_out[841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.265 0.070 622.335 ;
    END
  END rd_out[841]
  PIN rd_out[842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.405 0.070 622.475 ;
    END
  END rd_out[842]
  PIN rd_out[843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.545 0.070 622.615 ;
    END
  END rd_out[843]
  PIN rd_out[844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.685 0.070 622.755 ;
    END
  END rd_out[844]
  PIN rd_out[845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.825 0.070 622.895 ;
    END
  END rd_out[845]
  PIN rd_out[846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 622.965 0.070 623.035 ;
    END
  END rd_out[846]
  PIN rd_out[847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.105 0.070 623.175 ;
    END
  END rd_out[847]
  PIN rd_out[848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.245 0.070 623.315 ;
    END
  END rd_out[848]
  PIN rd_out[849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.385 0.070 623.455 ;
    END
  END rd_out[849]
  PIN rd_out[850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.525 0.070 623.595 ;
    END
  END rd_out[850]
  PIN rd_out[851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.665 0.070 623.735 ;
    END
  END rd_out[851]
  PIN rd_out[852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.805 0.070 623.875 ;
    END
  END rd_out[852]
  PIN rd_out[853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 623.945 0.070 624.015 ;
    END
  END rd_out[853]
  PIN rd_out[854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.085 0.070 624.155 ;
    END
  END rd_out[854]
  PIN rd_out[855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.225 0.070 624.295 ;
    END
  END rd_out[855]
  PIN rd_out[856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.365 0.070 624.435 ;
    END
  END rd_out[856]
  PIN rd_out[857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.505 0.070 624.575 ;
    END
  END rd_out[857]
  PIN rd_out[858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.645 0.070 624.715 ;
    END
  END rd_out[858]
  PIN rd_out[859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.785 0.070 624.855 ;
    END
  END rd_out[859]
  PIN rd_out[860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 624.925 0.070 624.995 ;
    END
  END rd_out[860]
  PIN rd_out[861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.065 0.070 625.135 ;
    END
  END rd_out[861]
  PIN rd_out[862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.205 0.070 625.275 ;
    END
  END rd_out[862]
  PIN rd_out[863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.345 0.070 625.415 ;
    END
  END rd_out[863]
  PIN rd_out[864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.485 0.070 625.555 ;
    END
  END rd_out[864]
  PIN rd_out[865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.625 0.070 625.695 ;
    END
  END rd_out[865]
  PIN rd_out[866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.765 0.070 625.835 ;
    END
  END rd_out[866]
  PIN rd_out[867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 625.905 0.070 625.975 ;
    END
  END rd_out[867]
  PIN rd_out[868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.045 0.070 626.115 ;
    END
  END rd_out[868]
  PIN rd_out[869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.185 0.070 626.255 ;
    END
  END rd_out[869]
  PIN rd_out[870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.325 0.070 626.395 ;
    END
  END rd_out[870]
  PIN rd_out[871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.465 0.070 626.535 ;
    END
  END rd_out[871]
  PIN rd_out[872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.605 0.070 626.675 ;
    END
  END rd_out[872]
  PIN rd_out[873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.745 0.070 626.815 ;
    END
  END rd_out[873]
  PIN rd_out[874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 626.885 0.070 626.955 ;
    END
  END rd_out[874]
  PIN rd_out[875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.025 0.070 627.095 ;
    END
  END rd_out[875]
  PIN rd_out[876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.165 0.070 627.235 ;
    END
  END rd_out[876]
  PIN rd_out[877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.305 0.070 627.375 ;
    END
  END rd_out[877]
  PIN rd_out[878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.445 0.070 627.515 ;
    END
  END rd_out[878]
  PIN rd_out[879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.585 0.070 627.655 ;
    END
  END rd_out[879]
  PIN rd_out[880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.725 0.070 627.795 ;
    END
  END rd_out[880]
  PIN rd_out[881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 627.865 0.070 627.935 ;
    END
  END rd_out[881]
  PIN rd_out[882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.005 0.070 628.075 ;
    END
  END rd_out[882]
  PIN rd_out[883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.145 0.070 628.215 ;
    END
  END rd_out[883]
  PIN rd_out[884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.285 0.070 628.355 ;
    END
  END rd_out[884]
  PIN rd_out[885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.425 0.070 628.495 ;
    END
  END rd_out[885]
  PIN rd_out[886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.565 0.070 628.635 ;
    END
  END rd_out[886]
  PIN rd_out[887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.705 0.070 628.775 ;
    END
  END rd_out[887]
  PIN rd_out[888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.845 0.070 628.915 ;
    END
  END rd_out[888]
  PIN rd_out[889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 628.985 0.070 629.055 ;
    END
  END rd_out[889]
  PIN rd_out[890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.125 0.070 629.195 ;
    END
  END rd_out[890]
  PIN rd_out[891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.265 0.070 629.335 ;
    END
  END rd_out[891]
  PIN rd_out[892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.405 0.070 629.475 ;
    END
  END rd_out[892]
  PIN rd_out[893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.545 0.070 629.615 ;
    END
  END rd_out[893]
  PIN rd_out[894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.685 0.070 629.755 ;
    END
  END rd_out[894]
  PIN rd_out[895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.825 0.070 629.895 ;
    END
  END rd_out[895]
  PIN rd_out[896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 629.965 0.070 630.035 ;
    END
  END rd_out[896]
  PIN rd_out[897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.105 0.070 630.175 ;
    END
  END rd_out[897]
  PIN rd_out[898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.245 0.070 630.315 ;
    END
  END rd_out[898]
  PIN rd_out[899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.385 0.070 630.455 ;
    END
  END rd_out[899]
  PIN rd_out[900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.525 0.070 630.595 ;
    END
  END rd_out[900]
  PIN rd_out[901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.665 0.070 630.735 ;
    END
  END rd_out[901]
  PIN rd_out[902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.805 0.070 630.875 ;
    END
  END rd_out[902]
  PIN rd_out[903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 630.945 0.070 631.015 ;
    END
  END rd_out[903]
  PIN rd_out[904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.085 0.070 631.155 ;
    END
  END rd_out[904]
  PIN rd_out[905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.225 0.070 631.295 ;
    END
  END rd_out[905]
  PIN rd_out[906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.365 0.070 631.435 ;
    END
  END rd_out[906]
  PIN rd_out[907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.505 0.070 631.575 ;
    END
  END rd_out[907]
  PIN rd_out[908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.645 0.070 631.715 ;
    END
  END rd_out[908]
  PIN rd_out[909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.785 0.070 631.855 ;
    END
  END rd_out[909]
  PIN rd_out[910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 631.925 0.070 631.995 ;
    END
  END rd_out[910]
  PIN rd_out[911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.065 0.070 632.135 ;
    END
  END rd_out[911]
  PIN rd_out[912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.205 0.070 632.275 ;
    END
  END rd_out[912]
  PIN rd_out[913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.345 0.070 632.415 ;
    END
  END rd_out[913]
  PIN rd_out[914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.485 0.070 632.555 ;
    END
  END rd_out[914]
  PIN rd_out[915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.625 0.070 632.695 ;
    END
  END rd_out[915]
  PIN rd_out[916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.765 0.070 632.835 ;
    END
  END rd_out[916]
  PIN rd_out[917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 632.905 0.070 632.975 ;
    END
  END rd_out[917]
  PIN rd_out[918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.045 0.070 633.115 ;
    END
  END rd_out[918]
  PIN rd_out[919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.185 0.070 633.255 ;
    END
  END rd_out[919]
  PIN rd_out[920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.325 0.070 633.395 ;
    END
  END rd_out[920]
  PIN rd_out[921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.465 0.070 633.535 ;
    END
  END rd_out[921]
  PIN rd_out[922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.605 0.070 633.675 ;
    END
  END rd_out[922]
  PIN rd_out[923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.745 0.070 633.815 ;
    END
  END rd_out[923]
  PIN rd_out[924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 633.885 0.070 633.955 ;
    END
  END rd_out[924]
  PIN rd_out[925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.025 0.070 634.095 ;
    END
  END rd_out[925]
  PIN rd_out[926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.165 0.070 634.235 ;
    END
  END rd_out[926]
  PIN rd_out[927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.305 0.070 634.375 ;
    END
  END rd_out[927]
  PIN rd_out[928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.445 0.070 634.515 ;
    END
  END rd_out[928]
  PIN rd_out[929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.585 0.070 634.655 ;
    END
  END rd_out[929]
  PIN rd_out[930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.725 0.070 634.795 ;
    END
  END rd_out[930]
  PIN rd_out[931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 634.865 0.070 634.935 ;
    END
  END rd_out[931]
  PIN rd_out[932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.005 0.070 635.075 ;
    END
  END rd_out[932]
  PIN rd_out[933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.145 0.070 635.215 ;
    END
  END rd_out[933]
  PIN rd_out[934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.285 0.070 635.355 ;
    END
  END rd_out[934]
  PIN rd_out[935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.425 0.070 635.495 ;
    END
  END rd_out[935]
  PIN rd_out[936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.565 0.070 635.635 ;
    END
  END rd_out[936]
  PIN rd_out[937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.705 0.070 635.775 ;
    END
  END rd_out[937]
  PIN rd_out[938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.845 0.070 635.915 ;
    END
  END rd_out[938]
  PIN rd_out[939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 635.985 0.070 636.055 ;
    END
  END rd_out[939]
  PIN rd_out[940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.125 0.070 636.195 ;
    END
  END rd_out[940]
  PIN rd_out[941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.265 0.070 636.335 ;
    END
  END rd_out[941]
  PIN rd_out[942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.405 0.070 636.475 ;
    END
  END rd_out[942]
  PIN rd_out[943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.545 0.070 636.615 ;
    END
  END rd_out[943]
  PIN rd_out[944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.685 0.070 636.755 ;
    END
  END rd_out[944]
  PIN rd_out[945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.825 0.070 636.895 ;
    END
  END rd_out[945]
  PIN rd_out[946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 636.965 0.070 637.035 ;
    END
  END rd_out[946]
  PIN rd_out[947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.105 0.070 637.175 ;
    END
  END rd_out[947]
  PIN rd_out[948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.245 0.070 637.315 ;
    END
  END rd_out[948]
  PIN rd_out[949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.385 0.070 637.455 ;
    END
  END rd_out[949]
  PIN rd_out[950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.525 0.070 637.595 ;
    END
  END rd_out[950]
  PIN rd_out[951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.665 0.070 637.735 ;
    END
  END rd_out[951]
  PIN rd_out[952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.805 0.070 637.875 ;
    END
  END rd_out[952]
  PIN rd_out[953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 637.945 0.070 638.015 ;
    END
  END rd_out[953]
  PIN rd_out[954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.085 0.070 638.155 ;
    END
  END rd_out[954]
  PIN rd_out[955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.225 0.070 638.295 ;
    END
  END rd_out[955]
  PIN rd_out[956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.365 0.070 638.435 ;
    END
  END rd_out[956]
  PIN rd_out[957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.505 0.070 638.575 ;
    END
  END rd_out[957]
  PIN rd_out[958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.645 0.070 638.715 ;
    END
  END rd_out[958]
  PIN rd_out[959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.785 0.070 638.855 ;
    END
  END rd_out[959]
  PIN rd_out[960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 638.925 0.070 638.995 ;
    END
  END rd_out[960]
  PIN rd_out[961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.065 0.070 639.135 ;
    END
  END rd_out[961]
  PIN rd_out[962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.205 0.070 639.275 ;
    END
  END rd_out[962]
  PIN rd_out[963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.345 0.070 639.415 ;
    END
  END rd_out[963]
  PIN rd_out[964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.485 0.070 639.555 ;
    END
  END rd_out[964]
  PIN rd_out[965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.625 0.070 639.695 ;
    END
  END rd_out[965]
  PIN rd_out[966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.765 0.070 639.835 ;
    END
  END rd_out[966]
  PIN rd_out[967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 639.905 0.070 639.975 ;
    END
  END rd_out[967]
  PIN rd_out[968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.045 0.070 640.115 ;
    END
  END rd_out[968]
  PIN rd_out[969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.185 0.070 640.255 ;
    END
  END rd_out[969]
  PIN rd_out[970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.325 0.070 640.395 ;
    END
  END rd_out[970]
  PIN rd_out[971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.465 0.070 640.535 ;
    END
  END rd_out[971]
  PIN rd_out[972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.605 0.070 640.675 ;
    END
  END rd_out[972]
  PIN rd_out[973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.745 0.070 640.815 ;
    END
  END rd_out[973]
  PIN rd_out[974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 640.885 0.070 640.955 ;
    END
  END rd_out[974]
  PIN rd_out[975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.025 0.070 641.095 ;
    END
  END rd_out[975]
  PIN rd_out[976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.165 0.070 641.235 ;
    END
  END rd_out[976]
  PIN rd_out[977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.305 0.070 641.375 ;
    END
  END rd_out[977]
  PIN rd_out[978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.445 0.070 641.515 ;
    END
  END rd_out[978]
  PIN rd_out[979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.585 0.070 641.655 ;
    END
  END rd_out[979]
  PIN rd_out[980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.725 0.070 641.795 ;
    END
  END rd_out[980]
  PIN rd_out[981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 641.865 0.070 641.935 ;
    END
  END rd_out[981]
  PIN rd_out[982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.005 0.070 642.075 ;
    END
  END rd_out[982]
  PIN rd_out[983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.145 0.070 642.215 ;
    END
  END rd_out[983]
  PIN rd_out[984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.285 0.070 642.355 ;
    END
  END rd_out[984]
  PIN rd_out[985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.425 0.070 642.495 ;
    END
  END rd_out[985]
  PIN rd_out[986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.565 0.070 642.635 ;
    END
  END rd_out[986]
  PIN rd_out[987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.705 0.070 642.775 ;
    END
  END rd_out[987]
  PIN rd_out[988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.845 0.070 642.915 ;
    END
  END rd_out[988]
  PIN rd_out[989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 642.985 0.070 643.055 ;
    END
  END rd_out[989]
  PIN rd_out[990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.125 0.070 643.195 ;
    END
  END rd_out[990]
  PIN rd_out[991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.265 0.070 643.335 ;
    END
  END rd_out[991]
  PIN rd_out[992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.405 0.070 643.475 ;
    END
  END rd_out[992]
  PIN rd_out[993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.545 0.070 643.615 ;
    END
  END rd_out[993]
  PIN rd_out[994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.685 0.070 643.755 ;
    END
  END rd_out[994]
  PIN rd_out[995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.825 0.070 643.895 ;
    END
  END rd_out[995]
  PIN rd_out[996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 643.965 0.070 644.035 ;
    END
  END rd_out[996]
  PIN rd_out[997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.105 0.070 644.175 ;
    END
  END rd_out[997]
  PIN rd_out[998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.245 0.070 644.315 ;
    END
  END rd_out[998]
  PIN rd_out[999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.385 0.070 644.455 ;
    END
  END rd_out[999]
  PIN rd_out[1000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.525 0.070 644.595 ;
    END
  END rd_out[1000]
  PIN rd_out[1001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.665 0.070 644.735 ;
    END
  END rd_out[1001]
  PIN rd_out[1002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.805 0.070 644.875 ;
    END
  END rd_out[1002]
  PIN rd_out[1003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 644.945 0.070 645.015 ;
    END
  END rd_out[1003]
  PIN rd_out[1004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.085 0.070 645.155 ;
    END
  END rd_out[1004]
  PIN rd_out[1005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.225 0.070 645.295 ;
    END
  END rd_out[1005]
  PIN rd_out[1006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.365 0.070 645.435 ;
    END
  END rd_out[1006]
  PIN rd_out[1007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.505 0.070 645.575 ;
    END
  END rd_out[1007]
  PIN rd_out[1008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.645 0.070 645.715 ;
    END
  END rd_out[1008]
  PIN rd_out[1009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.785 0.070 645.855 ;
    END
  END rd_out[1009]
  PIN rd_out[1010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 645.925 0.070 645.995 ;
    END
  END rd_out[1010]
  PIN rd_out[1011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.065 0.070 646.135 ;
    END
  END rd_out[1011]
  PIN rd_out[1012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.205 0.070 646.275 ;
    END
  END rd_out[1012]
  PIN rd_out[1013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.345 0.070 646.415 ;
    END
  END rd_out[1013]
  PIN rd_out[1014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.485 0.070 646.555 ;
    END
  END rd_out[1014]
  PIN rd_out[1015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.625 0.070 646.695 ;
    END
  END rd_out[1015]
  PIN rd_out[1016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.765 0.070 646.835 ;
    END
  END rd_out[1016]
  PIN rd_out[1017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 646.905 0.070 646.975 ;
    END
  END rd_out[1017]
  PIN rd_out[1018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.045 0.070 647.115 ;
    END
  END rd_out[1018]
  PIN rd_out[1019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.185 0.070 647.255 ;
    END
  END rd_out[1019]
  PIN rd_out[1020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.325 0.070 647.395 ;
    END
  END rd_out[1020]
  PIN rd_out[1021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.465 0.070 647.535 ;
    END
  END rd_out[1021]
  PIN rd_out[1022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.605 0.070 647.675 ;
    END
  END rd_out[1022]
  PIN rd_out[1023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.745 0.070 647.815 ;
    END
  END rd_out[1023]
  PIN rd_out[1024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 647.885 0.070 647.955 ;
    END
  END rd_out[1024]
  PIN rd_out[1025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.025 0.070 648.095 ;
    END
  END rd_out[1025]
  PIN rd_out[1026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.165 0.070 648.235 ;
    END
  END rd_out[1026]
  PIN rd_out[1027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.305 0.070 648.375 ;
    END
  END rd_out[1027]
  PIN rd_out[1028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.445 0.070 648.515 ;
    END
  END rd_out[1028]
  PIN rd_out[1029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.585 0.070 648.655 ;
    END
  END rd_out[1029]
  PIN rd_out[1030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.725 0.070 648.795 ;
    END
  END rd_out[1030]
  PIN rd_out[1031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 648.865 0.070 648.935 ;
    END
  END rd_out[1031]
  PIN rd_out[1032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.005 0.070 649.075 ;
    END
  END rd_out[1032]
  PIN rd_out[1033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.145 0.070 649.215 ;
    END
  END rd_out[1033]
  PIN rd_out[1034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.285 0.070 649.355 ;
    END
  END rd_out[1034]
  PIN rd_out[1035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.425 0.070 649.495 ;
    END
  END rd_out[1035]
  PIN rd_out[1036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.565 0.070 649.635 ;
    END
  END rd_out[1036]
  PIN rd_out[1037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.705 0.070 649.775 ;
    END
  END rd_out[1037]
  PIN rd_out[1038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.845 0.070 649.915 ;
    END
  END rd_out[1038]
  PIN rd_out[1039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 649.985 0.070 650.055 ;
    END
  END rd_out[1039]
  PIN rd_out[1040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.125 0.070 650.195 ;
    END
  END rd_out[1040]
  PIN rd_out[1041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.265 0.070 650.335 ;
    END
  END rd_out[1041]
  PIN rd_out[1042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.405 0.070 650.475 ;
    END
  END rd_out[1042]
  PIN rd_out[1043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.545 0.070 650.615 ;
    END
  END rd_out[1043]
  PIN rd_out[1044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.685 0.070 650.755 ;
    END
  END rd_out[1044]
  PIN rd_out[1045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.825 0.070 650.895 ;
    END
  END rd_out[1045]
  PIN rd_out[1046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 650.965 0.070 651.035 ;
    END
  END rd_out[1046]
  PIN rd_out[1047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.105 0.070 651.175 ;
    END
  END rd_out[1047]
  PIN rd_out[1048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.245 0.070 651.315 ;
    END
  END rd_out[1048]
  PIN rd_out[1049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.385 0.070 651.455 ;
    END
  END rd_out[1049]
  PIN rd_out[1050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.525 0.070 651.595 ;
    END
  END rd_out[1050]
  PIN rd_out[1051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.665 0.070 651.735 ;
    END
  END rd_out[1051]
  PIN rd_out[1052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.805 0.070 651.875 ;
    END
  END rd_out[1052]
  PIN rd_out[1053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 651.945 0.070 652.015 ;
    END
  END rd_out[1053]
  PIN rd_out[1054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.085 0.070 652.155 ;
    END
  END rd_out[1054]
  PIN rd_out[1055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.225 0.070 652.295 ;
    END
  END rd_out[1055]
  PIN rd_out[1056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.365 0.070 652.435 ;
    END
  END rd_out[1056]
  PIN rd_out[1057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.505 0.070 652.575 ;
    END
  END rd_out[1057]
  PIN rd_out[1058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.645 0.070 652.715 ;
    END
  END rd_out[1058]
  PIN rd_out[1059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.785 0.070 652.855 ;
    END
  END rd_out[1059]
  PIN rd_out[1060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 652.925 0.070 652.995 ;
    END
  END rd_out[1060]
  PIN rd_out[1061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.065 0.070 653.135 ;
    END
  END rd_out[1061]
  PIN rd_out[1062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.205 0.070 653.275 ;
    END
  END rd_out[1062]
  PIN rd_out[1063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.345 0.070 653.415 ;
    END
  END rd_out[1063]
  PIN rd_out[1064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.485 0.070 653.555 ;
    END
  END rd_out[1064]
  PIN rd_out[1065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.625 0.070 653.695 ;
    END
  END rd_out[1065]
  PIN rd_out[1066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.765 0.070 653.835 ;
    END
  END rd_out[1066]
  PIN rd_out[1067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 653.905 0.070 653.975 ;
    END
  END rd_out[1067]
  PIN rd_out[1068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.045 0.070 654.115 ;
    END
  END rd_out[1068]
  PIN rd_out[1069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.185 0.070 654.255 ;
    END
  END rd_out[1069]
  PIN rd_out[1070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.325 0.070 654.395 ;
    END
  END rd_out[1070]
  PIN rd_out[1071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.465 0.070 654.535 ;
    END
  END rd_out[1071]
  PIN rd_out[1072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.605 0.070 654.675 ;
    END
  END rd_out[1072]
  PIN rd_out[1073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.745 0.070 654.815 ;
    END
  END rd_out[1073]
  PIN rd_out[1074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 654.885 0.070 654.955 ;
    END
  END rd_out[1074]
  PIN rd_out[1075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.025 0.070 655.095 ;
    END
  END rd_out[1075]
  PIN rd_out[1076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.165 0.070 655.235 ;
    END
  END rd_out[1076]
  PIN rd_out[1077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.305 0.070 655.375 ;
    END
  END rd_out[1077]
  PIN rd_out[1078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.445 0.070 655.515 ;
    END
  END rd_out[1078]
  PIN rd_out[1079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.585 0.070 655.655 ;
    END
  END rd_out[1079]
  PIN rd_out[1080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.725 0.070 655.795 ;
    END
  END rd_out[1080]
  PIN rd_out[1081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 655.865 0.070 655.935 ;
    END
  END rd_out[1081]
  PIN rd_out[1082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.005 0.070 656.075 ;
    END
  END rd_out[1082]
  PIN rd_out[1083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.145 0.070 656.215 ;
    END
  END rd_out[1083]
  PIN rd_out[1084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.285 0.070 656.355 ;
    END
  END rd_out[1084]
  PIN rd_out[1085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.425 0.070 656.495 ;
    END
  END rd_out[1085]
  PIN rd_out[1086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.565 0.070 656.635 ;
    END
  END rd_out[1086]
  PIN rd_out[1087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.705 0.070 656.775 ;
    END
  END rd_out[1087]
  PIN rd_out[1088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.845 0.070 656.915 ;
    END
  END rd_out[1088]
  PIN rd_out[1089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 656.985 0.070 657.055 ;
    END
  END rd_out[1089]
  PIN rd_out[1090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.125 0.070 657.195 ;
    END
  END rd_out[1090]
  PIN rd_out[1091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.265 0.070 657.335 ;
    END
  END rd_out[1091]
  PIN rd_out[1092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.405 0.070 657.475 ;
    END
  END rd_out[1092]
  PIN rd_out[1093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.545 0.070 657.615 ;
    END
  END rd_out[1093]
  PIN rd_out[1094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.685 0.070 657.755 ;
    END
  END rd_out[1094]
  PIN rd_out[1095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.825 0.070 657.895 ;
    END
  END rd_out[1095]
  PIN rd_out[1096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 657.965 0.070 658.035 ;
    END
  END rd_out[1096]
  PIN rd_out[1097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.105 0.070 658.175 ;
    END
  END rd_out[1097]
  PIN rd_out[1098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.245 0.070 658.315 ;
    END
  END rd_out[1098]
  PIN rd_out[1099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.385 0.070 658.455 ;
    END
  END rd_out[1099]
  PIN rd_out[1100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.525 0.070 658.595 ;
    END
  END rd_out[1100]
  PIN rd_out[1101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.665 0.070 658.735 ;
    END
  END rd_out[1101]
  PIN rd_out[1102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.805 0.070 658.875 ;
    END
  END rd_out[1102]
  PIN rd_out[1103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 658.945 0.070 659.015 ;
    END
  END rd_out[1103]
  PIN rd_out[1104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.085 0.070 659.155 ;
    END
  END rd_out[1104]
  PIN rd_out[1105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.225 0.070 659.295 ;
    END
  END rd_out[1105]
  PIN rd_out[1106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.365 0.070 659.435 ;
    END
  END rd_out[1106]
  PIN rd_out[1107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.505 0.070 659.575 ;
    END
  END rd_out[1107]
  PIN rd_out[1108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.645 0.070 659.715 ;
    END
  END rd_out[1108]
  PIN rd_out[1109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.785 0.070 659.855 ;
    END
  END rd_out[1109]
  PIN rd_out[1110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 659.925 0.070 659.995 ;
    END
  END rd_out[1110]
  PIN rd_out[1111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.065 0.070 660.135 ;
    END
  END rd_out[1111]
  PIN rd_out[1112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.205 0.070 660.275 ;
    END
  END rd_out[1112]
  PIN rd_out[1113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.345 0.070 660.415 ;
    END
  END rd_out[1113]
  PIN rd_out[1114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.485 0.070 660.555 ;
    END
  END rd_out[1114]
  PIN rd_out[1115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.625 0.070 660.695 ;
    END
  END rd_out[1115]
  PIN rd_out[1116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.765 0.070 660.835 ;
    END
  END rd_out[1116]
  PIN rd_out[1117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 660.905 0.070 660.975 ;
    END
  END rd_out[1117]
  PIN rd_out[1118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.045 0.070 661.115 ;
    END
  END rd_out[1118]
  PIN rd_out[1119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.185 0.070 661.255 ;
    END
  END rd_out[1119]
  PIN rd_out[1120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.325 0.070 661.395 ;
    END
  END rd_out[1120]
  PIN rd_out[1121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.465 0.070 661.535 ;
    END
  END rd_out[1121]
  PIN rd_out[1122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.605 0.070 661.675 ;
    END
  END rd_out[1122]
  PIN rd_out[1123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.745 0.070 661.815 ;
    END
  END rd_out[1123]
  PIN rd_out[1124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 661.885 0.070 661.955 ;
    END
  END rd_out[1124]
  PIN rd_out[1125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.025 0.070 662.095 ;
    END
  END rd_out[1125]
  PIN rd_out[1126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.165 0.070 662.235 ;
    END
  END rd_out[1126]
  PIN rd_out[1127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.305 0.070 662.375 ;
    END
  END rd_out[1127]
  PIN rd_out[1128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.445 0.070 662.515 ;
    END
  END rd_out[1128]
  PIN rd_out[1129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.585 0.070 662.655 ;
    END
  END rd_out[1129]
  PIN rd_out[1130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.725 0.070 662.795 ;
    END
  END rd_out[1130]
  PIN rd_out[1131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 662.865 0.070 662.935 ;
    END
  END rd_out[1131]
  PIN rd_out[1132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.005 0.070 663.075 ;
    END
  END rd_out[1132]
  PIN rd_out[1133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.145 0.070 663.215 ;
    END
  END rd_out[1133]
  PIN rd_out[1134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.285 0.070 663.355 ;
    END
  END rd_out[1134]
  PIN rd_out[1135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.425 0.070 663.495 ;
    END
  END rd_out[1135]
  PIN rd_out[1136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.565 0.070 663.635 ;
    END
  END rd_out[1136]
  PIN rd_out[1137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.705 0.070 663.775 ;
    END
  END rd_out[1137]
  PIN rd_out[1138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.845 0.070 663.915 ;
    END
  END rd_out[1138]
  PIN rd_out[1139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 663.985 0.070 664.055 ;
    END
  END rd_out[1139]
  PIN rd_out[1140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.125 0.070 664.195 ;
    END
  END rd_out[1140]
  PIN rd_out[1141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.265 0.070 664.335 ;
    END
  END rd_out[1141]
  PIN rd_out[1142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.405 0.070 664.475 ;
    END
  END rd_out[1142]
  PIN rd_out[1143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.545 0.070 664.615 ;
    END
  END rd_out[1143]
  PIN rd_out[1144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.685 0.070 664.755 ;
    END
  END rd_out[1144]
  PIN rd_out[1145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.825 0.070 664.895 ;
    END
  END rd_out[1145]
  PIN rd_out[1146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 664.965 0.070 665.035 ;
    END
  END rd_out[1146]
  PIN rd_out[1147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.105 0.070 665.175 ;
    END
  END rd_out[1147]
  PIN rd_out[1148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.245 0.070 665.315 ;
    END
  END rd_out[1148]
  PIN rd_out[1149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.385 0.070 665.455 ;
    END
  END rd_out[1149]
  PIN rd_out[1150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.525 0.070 665.595 ;
    END
  END rd_out[1150]
  PIN rd_out[1151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.665 0.070 665.735 ;
    END
  END rd_out[1151]
  PIN rd_out[1152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.805 0.070 665.875 ;
    END
  END rd_out[1152]
  PIN rd_out[1153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 665.945 0.070 666.015 ;
    END
  END rd_out[1153]
  PIN rd_out[1154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.085 0.070 666.155 ;
    END
  END rd_out[1154]
  PIN rd_out[1155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.225 0.070 666.295 ;
    END
  END rd_out[1155]
  PIN rd_out[1156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.365 0.070 666.435 ;
    END
  END rd_out[1156]
  PIN rd_out[1157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.505 0.070 666.575 ;
    END
  END rd_out[1157]
  PIN rd_out[1158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.645 0.070 666.715 ;
    END
  END rd_out[1158]
  PIN rd_out[1159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.785 0.070 666.855 ;
    END
  END rd_out[1159]
  PIN rd_out[1160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 666.925 0.070 666.995 ;
    END
  END rd_out[1160]
  PIN rd_out[1161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.065 0.070 667.135 ;
    END
  END rd_out[1161]
  PIN rd_out[1162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.205 0.070 667.275 ;
    END
  END rd_out[1162]
  PIN rd_out[1163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.345 0.070 667.415 ;
    END
  END rd_out[1163]
  PIN rd_out[1164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.485 0.070 667.555 ;
    END
  END rd_out[1164]
  PIN rd_out[1165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.625 0.070 667.695 ;
    END
  END rd_out[1165]
  PIN rd_out[1166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.765 0.070 667.835 ;
    END
  END rd_out[1166]
  PIN rd_out[1167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 667.905 0.070 667.975 ;
    END
  END rd_out[1167]
  PIN rd_out[1168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.045 0.070 668.115 ;
    END
  END rd_out[1168]
  PIN rd_out[1169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.185 0.070 668.255 ;
    END
  END rd_out[1169]
  PIN rd_out[1170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.325 0.070 668.395 ;
    END
  END rd_out[1170]
  PIN rd_out[1171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.465 0.070 668.535 ;
    END
  END rd_out[1171]
  PIN rd_out[1172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.605 0.070 668.675 ;
    END
  END rd_out[1172]
  PIN rd_out[1173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.745 0.070 668.815 ;
    END
  END rd_out[1173]
  PIN rd_out[1174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 668.885 0.070 668.955 ;
    END
  END rd_out[1174]
  PIN rd_out[1175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.025 0.070 669.095 ;
    END
  END rd_out[1175]
  PIN rd_out[1176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.165 0.070 669.235 ;
    END
  END rd_out[1176]
  PIN rd_out[1177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.305 0.070 669.375 ;
    END
  END rd_out[1177]
  PIN rd_out[1178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.445 0.070 669.515 ;
    END
  END rd_out[1178]
  PIN rd_out[1179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.585 0.070 669.655 ;
    END
  END rd_out[1179]
  PIN rd_out[1180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.725 0.070 669.795 ;
    END
  END rd_out[1180]
  PIN rd_out[1181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 669.865 0.070 669.935 ;
    END
  END rd_out[1181]
  PIN rd_out[1182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.005 0.070 670.075 ;
    END
  END rd_out[1182]
  PIN rd_out[1183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.145 0.070 670.215 ;
    END
  END rd_out[1183]
  PIN rd_out[1184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.285 0.070 670.355 ;
    END
  END rd_out[1184]
  PIN rd_out[1185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.425 0.070 670.495 ;
    END
  END rd_out[1185]
  PIN rd_out[1186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.565 0.070 670.635 ;
    END
  END rd_out[1186]
  PIN rd_out[1187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.705 0.070 670.775 ;
    END
  END rd_out[1187]
  PIN rd_out[1188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.845 0.070 670.915 ;
    END
  END rd_out[1188]
  PIN rd_out[1189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 670.985 0.070 671.055 ;
    END
  END rd_out[1189]
  PIN rd_out[1190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.125 0.070 671.195 ;
    END
  END rd_out[1190]
  PIN rd_out[1191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.265 0.070 671.335 ;
    END
  END rd_out[1191]
  PIN rd_out[1192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.405 0.070 671.475 ;
    END
  END rd_out[1192]
  PIN rd_out[1193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.545 0.070 671.615 ;
    END
  END rd_out[1193]
  PIN rd_out[1194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.685 0.070 671.755 ;
    END
  END rd_out[1194]
  PIN rd_out[1195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.825 0.070 671.895 ;
    END
  END rd_out[1195]
  PIN rd_out[1196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 671.965 0.070 672.035 ;
    END
  END rd_out[1196]
  PIN rd_out[1197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.105 0.070 672.175 ;
    END
  END rd_out[1197]
  PIN rd_out[1198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.245 0.070 672.315 ;
    END
  END rd_out[1198]
  PIN rd_out[1199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.385 0.070 672.455 ;
    END
  END rd_out[1199]
  PIN rd_out[1200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.525 0.070 672.595 ;
    END
  END rd_out[1200]
  PIN rd_out[1201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.665 0.070 672.735 ;
    END
  END rd_out[1201]
  PIN rd_out[1202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.805 0.070 672.875 ;
    END
  END rd_out[1202]
  PIN rd_out[1203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 672.945 0.070 673.015 ;
    END
  END rd_out[1203]
  PIN rd_out[1204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.085 0.070 673.155 ;
    END
  END rd_out[1204]
  PIN rd_out[1205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.225 0.070 673.295 ;
    END
  END rd_out[1205]
  PIN rd_out[1206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.365 0.070 673.435 ;
    END
  END rd_out[1206]
  PIN rd_out[1207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.505 0.070 673.575 ;
    END
  END rd_out[1207]
  PIN rd_out[1208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.645 0.070 673.715 ;
    END
  END rd_out[1208]
  PIN rd_out[1209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.785 0.070 673.855 ;
    END
  END rd_out[1209]
  PIN rd_out[1210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 673.925 0.070 673.995 ;
    END
  END rd_out[1210]
  PIN rd_out[1211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.065 0.070 674.135 ;
    END
  END rd_out[1211]
  PIN rd_out[1212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.205 0.070 674.275 ;
    END
  END rd_out[1212]
  PIN rd_out[1213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.345 0.070 674.415 ;
    END
  END rd_out[1213]
  PIN rd_out[1214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.485 0.070 674.555 ;
    END
  END rd_out[1214]
  PIN rd_out[1215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.625 0.070 674.695 ;
    END
  END rd_out[1215]
  PIN rd_out[1216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.765 0.070 674.835 ;
    END
  END rd_out[1216]
  PIN rd_out[1217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 674.905 0.070 674.975 ;
    END
  END rd_out[1217]
  PIN rd_out[1218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.045 0.070 675.115 ;
    END
  END rd_out[1218]
  PIN rd_out[1219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.185 0.070 675.255 ;
    END
  END rd_out[1219]
  PIN rd_out[1220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.325 0.070 675.395 ;
    END
  END rd_out[1220]
  PIN rd_out[1221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.465 0.070 675.535 ;
    END
  END rd_out[1221]
  PIN rd_out[1222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.605 0.070 675.675 ;
    END
  END rd_out[1222]
  PIN rd_out[1223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.745 0.070 675.815 ;
    END
  END rd_out[1223]
  PIN rd_out[1224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 675.885 0.070 675.955 ;
    END
  END rd_out[1224]
  PIN rd_out[1225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.025 0.070 676.095 ;
    END
  END rd_out[1225]
  PIN rd_out[1226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.165 0.070 676.235 ;
    END
  END rd_out[1226]
  PIN rd_out[1227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.305 0.070 676.375 ;
    END
  END rd_out[1227]
  PIN rd_out[1228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.445 0.070 676.515 ;
    END
  END rd_out[1228]
  PIN rd_out[1229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.585 0.070 676.655 ;
    END
  END rd_out[1229]
  PIN rd_out[1230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.725 0.070 676.795 ;
    END
  END rd_out[1230]
  PIN rd_out[1231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 676.865 0.070 676.935 ;
    END
  END rd_out[1231]
  PIN rd_out[1232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.005 0.070 677.075 ;
    END
  END rd_out[1232]
  PIN rd_out[1233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.145 0.070 677.215 ;
    END
  END rd_out[1233]
  PIN rd_out[1234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.285 0.070 677.355 ;
    END
  END rd_out[1234]
  PIN rd_out[1235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.425 0.070 677.495 ;
    END
  END rd_out[1235]
  PIN rd_out[1236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.565 0.070 677.635 ;
    END
  END rd_out[1236]
  PIN rd_out[1237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.705 0.070 677.775 ;
    END
  END rd_out[1237]
  PIN rd_out[1238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.845 0.070 677.915 ;
    END
  END rd_out[1238]
  PIN rd_out[1239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 677.985 0.070 678.055 ;
    END
  END rd_out[1239]
  PIN rd_out[1240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.125 0.070 678.195 ;
    END
  END rd_out[1240]
  PIN rd_out[1241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.265 0.070 678.335 ;
    END
  END rd_out[1241]
  PIN rd_out[1242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.405 0.070 678.475 ;
    END
  END rd_out[1242]
  PIN rd_out[1243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.545 0.070 678.615 ;
    END
  END rd_out[1243]
  PIN rd_out[1244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.685 0.070 678.755 ;
    END
  END rd_out[1244]
  PIN rd_out[1245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.825 0.070 678.895 ;
    END
  END rd_out[1245]
  PIN rd_out[1246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 678.965 0.070 679.035 ;
    END
  END rd_out[1246]
  PIN rd_out[1247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.105 0.070 679.175 ;
    END
  END rd_out[1247]
  PIN rd_out[1248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.245 0.070 679.315 ;
    END
  END rd_out[1248]
  PIN rd_out[1249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.385 0.070 679.455 ;
    END
  END rd_out[1249]
  PIN rd_out[1250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.525 0.070 679.595 ;
    END
  END rd_out[1250]
  PIN rd_out[1251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.665 0.070 679.735 ;
    END
  END rd_out[1251]
  PIN rd_out[1252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.805 0.070 679.875 ;
    END
  END rd_out[1252]
  PIN rd_out[1253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 679.945 0.070 680.015 ;
    END
  END rd_out[1253]
  PIN rd_out[1254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.085 0.070 680.155 ;
    END
  END rd_out[1254]
  PIN rd_out[1255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.225 0.070 680.295 ;
    END
  END rd_out[1255]
  PIN rd_out[1256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.365 0.070 680.435 ;
    END
  END rd_out[1256]
  PIN rd_out[1257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.505 0.070 680.575 ;
    END
  END rd_out[1257]
  PIN rd_out[1258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.645 0.070 680.715 ;
    END
  END rd_out[1258]
  PIN rd_out[1259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.785 0.070 680.855 ;
    END
  END rd_out[1259]
  PIN rd_out[1260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 680.925 0.070 680.995 ;
    END
  END rd_out[1260]
  PIN rd_out[1261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.065 0.070 681.135 ;
    END
  END rd_out[1261]
  PIN rd_out[1262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.205 0.070 681.275 ;
    END
  END rd_out[1262]
  PIN rd_out[1263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.345 0.070 681.415 ;
    END
  END rd_out[1263]
  PIN rd_out[1264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.485 0.070 681.555 ;
    END
  END rd_out[1264]
  PIN rd_out[1265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.625 0.070 681.695 ;
    END
  END rd_out[1265]
  PIN rd_out[1266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.765 0.070 681.835 ;
    END
  END rd_out[1266]
  PIN rd_out[1267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 681.905 0.070 681.975 ;
    END
  END rd_out[1267]
  PIN rd_out[1268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.045 0.070 682.115 ;
    END
  END rd_out[1268]
  PIN rd_out[1269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.185 0.070 682.255 ;
    END
  END rd_out[1269]
  PIN rd_out[1270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.325 0.070 682.395 ;
    END
  END rd_out[1270]
  PIN rd_out[1271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.465 0.070 682.535 ;
    END
  END rd_out[1271]
  PIN rd_out[1272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.605 0.070 682.675 ;
    END
  END rd_out[1272]
  PIN rd_out[1273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.745 0.070 682.815 ;
    END
  END rd_out[1273]
  PIN rd_out[1274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 682.885 0.070 682.955 ;
    END
  END rd_out[1274]
  PIN rd_out[1275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.025 0.070 683.095 ;
    END
  END rd_out[1275]
  PIN rd_out[1276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.165 0.070 683.235 ;
    END
  END rd_out[1276]
  PIN rd_out[1277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.305 0.070 683.375 ;
    END
  END rd_out[1277]
  PIN rd_out[1278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.445 0.070 683.515 ;
    END
  END rd_out[1278]
  PIN rd_out[1279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.585 0.070 683.655 ;
    END
  END rd_out[1279]
  PIN rd_out[1280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.725 0.070 683.795 ;
    END
  END rd_out[1280]
  PIN rd_out[1281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 683.865 0.070 683.935 ;
    END
  END rd_out[1281]
  PIN rd_out[1282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.005 0.070 684.075 ;
    END
  END rd_out[1282]
  PIN rd_out[1283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.145 0.070 684.215 ;
    END
  END rd_out[1283]
  PIN rd_out[1284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.285 0.070 684.355 ;
    END
  END rd_out[1284]
  PIN rd_out[1285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.425 0.070 684.495 ;
    END
  END rd_out[1285]
  PIN rd_out[1286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.565 0.070 684.635 ;
    END
  END rd_out[1286]
  PIN rd_out[1287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.705 0.070 684.775 ;
    END
  END rd_out[1287]
  PIN rd_out[1288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.845 0.070 684.915 ;
    END
  END rd_out[1288]
  PIN rd_out[1289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 684.985 0.070 685.055 ;
    END
  END rd_out[1289]
  PIN rd_out[1290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.125 0.070 685.195 ;
    END
  END rd_out[1290]
  PIN rd_out[1291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.265 0.070 685.335 ;
    END
  END rd_out[1291]
  PIN rd_out[1292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.405 0.070 685.475 ;
    END
  END rd_out[1292]
  PIN rd_out[1293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.545 0.070 685.615 ;
    END
  END rd_out[1293]
  PIN rd_out[1294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.685 0.070 685.755 ;
    END
  END rd_out[1294]
  PIN rd_out[1295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.825 0.070 685.895 ;
    END
  END rd_out[1295]
  PIN rd_out[1296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 685.965 0.070 686.035 ;
    END
  END rd_out[1296]
  PIN rd_out[1297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.105 0.070 686.175 ;
    END
  END rd_out[1297]
  PIN rd_out[1298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.245 0.070 686.315 ;
    END
  END rd_out[1298]
  PIN rd_out[1299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.385 0.070 686.455 ;
    END
  END rd_out[1299]
  PIN rd_out[1300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.525 0.070 686.595 ;
    END
  END rd_out[1300]
  PIN rd_out[1301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.665 0.070 686.735 ;
    END
  END rd_out[1301]
  PIN rd_out[1302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.805 0.070 686.875 ;
    END
  END rd_out[1302]
  PIN rd_out[1303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 686.945 0.070 687.015 ;
    END
  END rd_out[1303]
  PIN rd_out[1304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.085 0.070 687.155 ;
    END
  END rd_out[1304]
  PIN rd_out[1305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.225 0.070 687.295 ;
    END
  END rd_out[1305]
  PIN rd_out[1306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.365 0.070 687.435 ;
    END
  END rd_out[1306]
  PIN rd_out[1307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.505 0.070 687.575 ;
    END
  END rd_out[1307]
  PIN rd_out[1308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.645 0.070 687.715 ;
    END
  END rd_out[1308]
  PIN rd_out[1309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.785 0.070 687.855 ;
    END
  END rd_out[1309]
  PIN rd_out[1310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 687.925 0.070 687.995 ;
    END
  END rd_out[1310]
  PIN rd_out[1311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.065 0.070 688.135 ;
    END
  END rd_out[1311]
  PIN rd_out[1312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.205 0.070 688.275 ;
    END
  END rd_out[1312]
  PIN rd_out[1313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.345 0.070 688.415 ;
    END
  END rd_out[1313]
  PIN rd_out[1314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.485 0.070 688.555 ;
    END
  END rd_out[1314]
  PIN rd_out[1315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.625 0.070 688.695 ;
    END
  END rd_out[1315]
  PIN rd_out[1316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.765 0.070 688.835 ;
    END
  END rd_out[1316]
  PIN rd_out[1317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 688.905 0.070 688.975 ;
    END
  END rd_out[1317]
  PIN rd_out[1318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.045 0.070 689.115 ;
    END
  END rd_out[1318]
  PIN rd_out[1319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.185 0.070 689.255 ;
    END
  END rd_out[1319]
  PIN rd_out[1320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.325 0.070 689.395 ;
    END
  END rd_out[1320]
  PIN rd_out[1321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.465 0.070 689.535 ;
    END
  END rd_out[1321]
  PIN rd_out[1322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.605 0.070 689.675 ;
    END
  END rd_out[1322]
  PIN rd_out[1323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.745 0.070 689.815 ;
    END
  END rd_out[1323]
  PIN rd_out[1324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 689.885 0.070 689.955 ;
    END
  END rd_out[1324]
  PIN rd_out[1325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.025 0.070 690.095 ;
    END
  END rd_out[1325]
  PIN rd_out[1326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.165 0.070 690.235 ;
    END
  END rd_out[1326]
  PIN rd_out[1327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.305 0.070 690.375 ;
    END
  END rd_out[1327]
  PIN rd_out[1328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.445 0.070 690.515 ;
    END
  END rd_out[1328]
  PIN rd_out[1329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.585 0.070 690.655 ;
    END
  END rd_out[1329]
  PIN rd_out[1330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.725 0.070 690.795 ;
    END
  END rd_out[1330]
  PIN rd_out[1331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 690.865 0.070 690.935 ;
    END
  END rd_out[1331]
  PIN rd_out[1332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.005 0.070 691.075 ;
    END
  END rd_out[1332]
  PIN rd_out[1333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.145 0.070 691.215 ;
    END
  END rd_out[1333]
  PIN rd_out[1334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.285 0.070 691.355 ;
    END
  END rd_out[1334]
  PIN rd_out[1335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.425 0.070 691.495 ;
    END
  END rd_out[1335]
  PIN rd_out[1336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.565 0.070 691.635 ;
    END
  END rd_out[1336]
  PIN rd_out[1337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.705 0.070 691.775 ;
    END
  END rd_out[1337]
  PIN rd_out[1338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.845 0.070 691.915 ;
    END
  END rd_out[1338]
  PIN rd_out[1339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 691.985 0.070 692.055 ;
    END
  END rd_out[1339]
  PIN rd_out[1340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.125 0.070 692.195 ;
    END
  END rd_out[1340]
  PIN rd_out[1341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.265 0.070 692.335 ;
    END
  END rd_out[1341]
  PIN rd_out[1342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.405 0.070 692.475 ;
    END
  END rd_out[1342]
  PIN rd_out[1343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.545 0.070 692.615 ;
    END
  END rd_out[1343]
  PIN rd_out[1344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.685 0.070 692.755 ;
    END
  END rd_out[1344]
  PIN rd_out[1345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.825 0.070 692.895 ;
    END
  END rd_out[1345]
  PIN rd_out[1346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 692.965 0.070 693.035 ;
    END
  END rd_out[1346]
  PIN rd_out[1347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.105 0.070 693.175 ;
    END
  END rd_out[1347]
  PIN rd_out[1348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.245 0.070 693.315 ;
    END
  END rd_out[1348]
  PIN rd_out[1349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.385 0.070 693.455 ;
    END
  END rd_out[1349]
  PIN rd_out[1350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.525 0.070 693.595 ;
    END
  END rd_out[1350]
  PIN rd_out[1351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.665 0.070 693.735 ;
    END
  END rd_out[1351]
  PIN rd_out[1352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.805 0.070 693.875 ;
    END
  END rd_out[1352]
  PIN rd_out[1353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 693.945 0.070 694.015 ;
    END
  END rd_out[1353]
  PIN rd_out[1354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.085 0.070 694.155 ;
    END
  END rd_out[1354]
  PIN rd_out[1355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.225 0.070 694.295 ;
    END
  END rd_out[1355]
  PIN rd_out[1356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.365 0.070 694.435 ;
    END
  END rd_out[1356]
  PIN rd_out[1357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.505 0.070 694.575 ;
    END
  END rd_out[1357]
  PIN rd_out[1358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.645 0.070 694.715 ;
    END
  END rd_out[1358]
  PIN rd_out[1359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.785 0.070 694.855 ;
    END
  END rd_out[1359]
  PIN rd_out[1360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 694.925 0.070 694.995 ;
    END
  END rd_out[1360]
  PIN rd_out[1361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.065 0.070 695.135 ;
    END
  END rd_out[1361]
  PIN rd_out[1362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.205 0.070 695.275 ;
    END
  END rd_out[1362]
  PIN rd_out[1363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.345 0.070 695.415 ;
    END
  END rd_out[1363]
  PIN rd_out[1364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.485 0.070 695.555 ;
    END
  END rd_out[1364]
  PIN rd_out[1365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.625 0.070 695.695 ;
    END
  END rd_out[1365]
  PIN rd_out[1366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.765 0.070 695.835 ;
    END
  END rd_out[1366]
  PIN rd_out[1367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 695.905 0.070 695.975 ;
    END
  END rd_out[1367]
  PIN rd_out[1368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.045 0.070 696.115 ;
    END
  END rd_out[1368]
  PIN rd_out[1369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.185 0.070 696.255 ;
    END
  END rd_out[1369]
  PIN rd_out[1370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.325 0.070 696.395 ;
    END
  END rd_out[1370]
  PIN rd_out[1371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.465 0.070 696.535 ;
    END
  END rd_out[1371]
  PIN rd_out[1372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.605 0.070 696.675 ;
    END
  END rd_out[1372]
  PIN rd_out[1373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.745 0.070 696.815 ;
    END
  END rd_out[1373]
  PIN rd_out[1374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 696.885 0.070 696.955 ;
    END
  END rd_out[1374]
  PIN rd_out[1375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.025 0.070 697.095 ;
    END
  END rd_out[1375]
  PIN rd_out[1376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.165 0.070 697.235 ;
    END
  END rd_out[1376]
  PIN rd_out[1377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.305 0.070 697.375 ;
    END
  END rd_out[1377]
  PIN rd_out[1378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.445 0.070 697.515 ;
    END
  END rd_out[1378]
  PIN rd_out[1379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.585 0.070 697.655 ;
    END
  END rd_out[1379]
  PIN rd_out[1380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.725 0.070 697.795 ;
    END
  END rd_out[1380]
  PIN rd_out[1381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 697.865 0.070 697.935 ;
    END
  END rd_out[1381]
  PIN rd_out[1382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.005 0.070 698.075 ;
    END
  END rd_out[1382]
  PIN rd_out[1383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.145 0.070 698.215 ;
    END
  END rd_out[1383]
  PIN rd_out[1384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.285 0.070 698.355 ;
    END
  END rd_out[1384]
  PIN rd_out[1385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.425 0.070 698.495 ;
    END
  END rd_out[1385]
  PIN rd_out[1386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.565 0.070 698.635 ;
    END
  END rd_out[1386]
  PIN rd_out[1387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.705 0.070 698.775 ;
    END
  END rd_out[1387]
  PIN rd_out[1388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.845 0.070 698.915 ;
    END
  END rd_out[1388]
  PIN rd_out[1389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 698.985 0.070 699.055 ;
    END
  END rd_out[1389]
  PIN rd_out[1390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.125 0.070 699.195 ;
    END
  END rd_out[1390]
  PIN rd_out[1391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.265 0.070 699.335 ;
    END
  END rd_out[1391]
  PIN rd_out[1392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.405 0.070 699.475 ;
    END
  END rd_out[1392]
  PIN rd_out[1393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.545 0.070 699.615 ;
    END
  END rd_out[1393]
  PIN rd_out[1394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.685 0.070 699.755 ;
    END
  END rd_out[1394]
  PIN rd_out[1395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.825 0.070 699.895 ;
    END
  END rd_out[1395]
  PIN rd_out[1396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 699.965 0.070 700.035 ;
    END
  END rd_out[1396]
  PIN rd_out[1397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.105 0.070 700.175 ;
    END
  END rd_out[1397]
  PIN rd_out[1398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.245 0.070 700.315 ;
    END
  END rd_out[1398]
  PIN rd_out[1399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.385 0.070 700.455 ;
    END
  END rd_out[1399]
  PIN rd_out[1400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.525 0.070 700.595 ;
    END
  END rd_out[1400]
  PIN rd_out[1401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.665 0.070 700.735 ;
    END
  END rd_out[1401]
  PIN rd_out[1402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.805 0.070 700.875 ;
    END
  END rd_out[1402]
  PIN rd_out[1403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 700.945 0.070 701.015 ;
    END
  END rd_out[1403]
  PIN rd_out[1404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.085 0.070 701.155 ;
    END
  END rd_out[1404]
  PIN rd_out[1405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.225 0.070 701.295 ;
    END
  END rd_out[1405]
  PIN rd_out[1406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.365 0.070 701.435 ;
    END
  END rd_out[1406]
  PIN rd_out[1407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.505 0.070 701.575 ;
    END
  END rd_out[1407]
  PIN rd_out[1408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.645 0.070 701.715 ;
    END
  END rd_out[1408]
  PIN rd_out[1409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.785 0.070 701.855 ;
    END
  END rd_out[1409]
  PIN rd_out[1410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 701.925 0.070 701.995 ;
    END
  END rd_out[1410]
  PIN rd_out[1411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.065 0.070 702.135 ;
    END
  END rd_out[1411]
  PIN rd_out[1412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.205 0.070 702.275 ;
    END
  END rd_out[1412]
  PIN rd_out[1413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.345 0.070 702.415 ;
    END
  END rd_out[1413]
  PIN rd_out[1414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.485 0.070 702.555 ;
    END
  END rd_out[1414]
  PIN rd_out[1415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.625 0.070 702.695 ;
    END
  END rd_out[1415]
  PIN rd_out[1416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.765 0.070 702.835 ;
    END
  END rd_out[1416]
  PIN rd_out[1417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 702.905 0.070 702.975 ;
    END
  END rd_out[1417]
  PIN rd_out[1418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.045 0.070 703.115 ;
    END
  END rd_out[1418]
  PIN rd_out[1419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.185 0.070 703.255 ;
    END
  END rd_out[1419]
  PIN rd_out[1420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.325 0.070 703.395 ;
    END
  END rd_out[1420]
  PIN rd_out[1421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.465 0.070 703.535 ;
    END
  END rd_out[1421]
  PIN rd_out[1422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.605 0.070 703.675 ;
    END
  END rd_out[1422]
  PIN rd_out[1423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.745 0.070 703.815 ;
    END
  END rd_out[1423]
  PIN rd_out[1424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 703.885 0.070 703.955 ;
    END
  END rd_out[1424]
  PIN rd_out[1425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.025 0.070 704.095 ;
    END
  END rd_out[1425]
  PIN rd_out[1426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.165 0.070 704.235 ;
    END
  END rd_out[1426]
  PIN rd_out[1427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.305 0.070 704.375 ;
    END
  END rd_out[1427]
  PIN rd_out[1428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.445 0.070 704.515 ;
    END
  END rd_out[1428]
  PIN rd_out[1429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.585 0.070 704.655 ;
    END
  END rd_out[1429]
  PIN rd_out[1430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.725 0.070 704.795 ;
    END
  END rd_out[1430]
  PIN rd_out[1431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 704.865 0.070 704.935 ;
    END
  END rd_out[1431]
  PIN rd_out[1432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.005 0.070 705.075 ;
    END
  END rd_out[1432]
  PIN rd_out[1433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.145 0.070 705.215 ;
    END
  END rd_out[1433]
  PIN rd_out[1434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.285 0.070 705.355 ;
    END
  END rd_out[1434]
  PIN rd_out[1435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.425 0.070 705.495 ;
    END
  END rd_out[1435]
  PIN rd_out[1436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.565 0.070 705.635 ;
    END
  END rd_out[1436]
  PIN rd_out[1437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.705 0.070 705.775 ;
    END
  END rd_out[1437]
  PIN rd_out[1438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.845 0.070 705.915 ;
    END
  END rd_out[1438]
  PIN rd_out[1439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 705.985 0.070 706.055 ;
    END
  END rd_out[1439]
  PIN rd_out[1440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.125 0.070 706.195 ;
    END
  END rd_out[1440]
  PIN rd_out[1441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.265 0.070 706.335 ;
    END
  END rd_out[1441]
  PIN rd_out[1442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.405 0.070 706.475 ;
    END
  END rd_out[1442]
  PIN rd_out[1443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.545 0.070 706.615 ;
    END
  END rd_out[1443]
  PIN rd_out[1444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.685 0.070 706.755 ;
    END
  END rd_out[1444]
  PIN rd_out[1445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.825 0.070 706.895 ;
    END
  END rd_out[1445]
  PIN rd_out[1446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 706.965 0.070 707.035 ;
    END
  END rd_out[1446]
  PIN rd_out[1447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.105 0.070 707.175 ;
    END
  END rd_out[1447]
  PIN rd_out[1448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.245 0.070 707.315 ;
    END
  END rd_out[1448]
  PIN rd_out[1449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.385 0.070 707.455 ;
    END
  END rd_out[1449]
  PIN rd_out[1450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.525 0.070 707.595 ;
    END
  END rd_out[1450]
  PIN rd_out[1451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.665 0.070 707.735 ;
    END
  END rd_out[1451]
  PIN rd_out[1452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.805 0.070 707.875 ;
    END
  END rd_out[1452]
  PIN rd_out[1453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 707.945 0.070 708.015 ;
    END
  END rd_out[1453]
  PIN rd_out[1454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.085 0.070 708.155 ;
    END
  END rd_out[1454]
  PIN rd_out[1455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.225 0.070 708.295 ;
    END
  END rd_out[1455]
  PIN rd_out[1456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.365 0.070 708.435 ;
    END
  END rd_out[1456]
  PIN rd_out[1457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.505 0.070 708.575 ;
    END
  END rd_out[1457]
  PIN rd_out[1458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.645 0.070 708.715 ;
    END
  END rd_out[1458]
  PIN rd_out[1459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.785 0.070 708.855 ;
    END
  END rd_out[1459]
  PIN rd_out[1460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 708.925 0.070 708.995 ;
    END
  END rd_out[1460]
  PIN rd_out[1461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.065 0.070 709.135 ;
    END
  END rd_out[1461]
  PIN rd_out[1462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.205 0.070 709.275 ;
    END
  END rd_out[1462]
  PIN rd_out[1463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.345 0.070 709.415 ;
    END
  END rd_out[1463]
  PIN rd_out[1464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.485 0.070 709.555 ;
    END
  END rd_out[1464]
  PIN rd_out[1465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.625 0.070 709.695 ;
    END
  END rd_out[1465]
  PIN rd_out[1466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.765 0.070 709.835 ;
    END
  END rd_out[1466]
  PIN rd_out[1467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 709.905 0.070 709.975 ;
    END
  END rd_out[1467]
  PIN rd_out[1468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.045 0.070 710.115 ;
    END
  END rd_out[1468]
  PIN rd_out[1469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.185 0.070 710.255 ;
    END
  END rd_out[1469]
  PIN rd_out[1470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.325 0.070 710.395 ;
    END
  END rd_out[1470]
  PIN rd_out[1471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.465 0.070 710.535 ;
    END
  END rd_out[1471]
  PIN rd_out[1472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.605 0.070 710.675 ;
    END
  END rd_out[1472]
  PIN rd_out[1473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.745 0.070 710.815 ;
    END
  END rd_out[1473]
  PIN rd_out[1474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 710.885 0.070 710.955 ;
    END
  END rd_out[1474]
  PIN rd_out[1475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.025 0.070 711.095 ;
    END
  END rd_out[1475]
  PIN rd_out[1476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.165 0.070 711.235 ;
    END
  END rd_out[1476]
  PIN rd_out[1477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.305 0.070 711.375 ;
    END
  END rd_out[1477]
  PIN rd_out[1478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.445 0.070 711.515 ;
    END
  END rd_out[1478]
  PIN rd_out[1479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.585 0.070 711.655 ;
    END
  END rd_out[1479]
  PIN rd_out[1480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.725 0.070 711.795 ;
    END
  END rd_out[1480]
  PIN rd_out[1481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 711.865 0.070 711.935 ;
    END
  END rd_out[1481]
  PIN rd_out[1482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.005 0.070 712.075 ;
    END
  END rd_out[1482]
  PIN rd_out[1483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.145 0.070 712.215 ;
    END
  END rd_out[1483]
  PIN rd_out[1484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.285 0.070 712.355 ;
    END
  END rd_out[1484]
  PIN rd_out[1485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.425 0.070 712.495 ;
    END
  END rd_out[1485]
  PIN rd_out[1486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.565 0.070 712.635 ;
    END
  END rd_out[1486]
  PIN rd_out[1487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.705 0.070 712.775 ;
    END
  END rd_out[1487]
  PIN rd_out[1488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.845 0.070 712.915 ;
    END
  END rd_out[1488]
  PIN rd_out[1489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 712.985 0.070 713.055 ;
    END
  END rd_out[1489]
  PIN rd_out[1490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.125 0.070 713.195 ;
    END
  END rd_out[1490]
  PIN rd_out[1491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.265 0.070 713.335 ;
    END
  END rd_out[1491]
  PIN rd_out[1492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.405 0.070 713.475 ;
    END
  END rd_out[1492]
  PIN rd_out[1493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.545 0.070 713.615 ;
    END
  END rd_out[1493]
  PIN rd_out[1494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.685 0.070 713.755 ;
    END
  END rd_out[1494]
  PIN rd_out[1495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.825 0.070 713.895 ;
    END
  END rd_out[1495]
  PIN rd_out[1496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 713.965 0.070 714.035 ;
    END
  END rd_out[1496]
  PIN rd_out[1497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.105 0.070 714.175 ;
    END
  END rd_out[1497]
  PIN rd_out[1498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.245 0.070 714.315 ;
    END
  END rd_out[1498]
  PIN rd_out[1499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.385 0.070 714.455 ;
    END
  END rd_out[1499]
  PIN rd_out[1500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.525 0.070 714.595 ;
    END
  END rd_out[1500]
  PIN rd_out[1501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.665 0.070 714.735 ;
    END
  END rd_out[1501]
  PIN rd_out[1502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.805 0.070 714.875 ;
    END
  END rd_out[1502]
  PIN rd_out[1503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 714.945 0.070 715.015 ;
    END
  END rd_out[1503]
  PIN rd_out[1504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.085 0.070 715.155 ;
    END
  END rd_out[1504]
  PIN rd_out[1505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.225 0.070 715.295 ;
    END
  END rd_out[1505]
  PIN rd_out[1506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.365 0.070 715.435 ;
    END
  END rd_out[1506]
  PIN rd_out[1507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.505 0.070 715.575 ;
    END
  END rd_out[1507]
  PIN rd_out[1508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.645 0.070 715.715 ;
    END
  END rd_out[1508]
  PIN rd_out[1509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.785 0.070 715.855 ;
    END
  END rd_out[1509]
  PIN rd_out[1510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 715.925 0.070 715.995 ;
    END
  END rd_out[1510]
  PIN rd_out[1511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.065 0.070 716.135 ;
    END
  END rd_out[1511]
  PIN rd_out[1512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.205 0.070 716.275 ;
    END
  END rd_out[1512]
  PIN rd_out[1513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.345 0.070 716.415 ;
    END
  END rd_out[1513]
  PIN rd_out[1514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.485 0.070 716.555 ;
    END
  END rd_out[1514]
  PIN rd_out[1515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.625 0.070 716.695 ;
    END
  END rd_out[1515]
  PIN rd_out[1516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.765 0.070 716.835 ;
    END
  END rd_out[1516]
  PIN rd_out[1517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 716.905 0.070 716.975 ;
    END
  END rd_out[1517]
  PIN rd_out[1518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.045 0.070 717.115 ;
    END
  END rd_out[1518]
  PIN rd_out[1519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.185 0.070 717.255 ;
    END
  END rd_out[1519]
  PIN rd_out[1520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.325 0.070 717.395 ;
    END
  END rd_out[1520]
  PIN rd_out[1521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.465 0.070 717.535 ;
    END
  END rd_out[1521]
  PIN rd_out[1522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.605 0.070 717.675 ;
    END
  END rd_out[1522]
  PIN rd_out[1523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.745 0.070 717.815 ;
    END
  END rd_out[1523]
  PIN rd_out[1524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 717.885 0.070 717.955 ;
    END
  END rd_out[1524]
  PIN rd_out[1525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.025 0.070 718.095 ;
    END
  END rd_out[1525]
  PIN rd_out[1526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.165 0.070 718.235 ;
    END
  END rd_out[1526]
  PIN rd_out[1527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.305 0.070 718.375 ;
    END
  END rd_out[1527]
  PIN rd_out[1528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.445 0.070 718.515 ;
    END
  END rd_out[1528]
  PIN rd_out[1529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.585 0.070 718.655 ;
    END
  END rd_out[1529]
  PIN rd_out[1530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.725 0.070 718.795 ;
    END
  END rd_out[1530]
  PIN rd_out[1531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 718.865 0.070 718.935 ;
    END
  END rd_out[1531]
  PIN rd_out[1532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.005 0.070 719.075 ;
    END
  END rd_out[1532]
  PIN rd_out[1533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.145 0.070 719.215 ;
    END
  END rd_out[1533]
  PIN rd_out[1534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.285 0.070 719.355 ;
    END
  END rd_out[1534]
  PIN rd_out[1535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.425 0.070 719.495 ;
    END
  END rd_out[1535]
  PIN rd_out[1536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.565 0.070 719.635 ;
    END
  END rd_out[1536]
  PIN rd_out[1537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.705 0.070 719.775 ;
    END
  END rd_out[1537]
  PIN rd_out[1538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.845 0.070 719.915 ;
    END
  END rd_out[1538]
  PIN rd_out[1539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 719.985 0.070 720.055 ;
    END
  END rd_out[1539]
  PIN rd_out[1540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.125 0.070 720.195 ;
    END
  END rd_out[1540]
  PIN rd_out[1541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.265 0.070 720.335 ;
    END
  END rd_out[1541]
  PIN rd_out[1542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.405 0.070 720.475 ;
    END
  END rd_out[1542]
  PIN rd_out[1543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.545 0.070 720.615 ;
    END
  END rd_out[1543]
  PIN rd_out[1544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.685 0.070 720.755 ;
    END
  END rd_out[1544]
  PIN rd_out[1545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.825 0.070 720.895 ;
    END
  END rd_out[1545]
  PIN rd_out[1546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 720.965 0.070 721.035 ;
    END
  END rd_out[1546]
  PIN rd_out[1547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.105 0.070 721.175 ;
    END
  END rd_out[1547]
  PIN rd_out[1548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.245 0.070 721.315 ;
    END
  END rd_out[1548]
  PIN rd_out[1549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.385 0.070 721.455 ;
    END
  END rd_out[1549]
  PIN rd_out[1550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.525 0.070 721.595 ;
    END
  END rd_out[1550]
  PIN rd_out[1551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.665 0.070 721.735 ;
    END
  END rd_out[1551]
  PIN rd_out[1552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.805 0.070 721.875 ;
    END
  END rd_out[1552]
  PIN rd_out[1553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 721.945 0.070 722.015 ;
    END
  END rd_out[1553]
  PIN rd_out[1554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.085 0.070 722.155 ;
    END
  END rd_out[1554]
  PIN rd_out[1555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.225 0.070 722.295 ;
    END
  END rd_out[1555]
  PIN rd_out[1556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.365 0.070 722.435 ;
    END
  END rd_out[1556]
  PIN rd_out[1557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.505 0.070 722.575 ;
    END
  END rd_out[1557]
  PIN rd_out[1558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.645 0.070 722.715 ;
    END
  END rd_out[1558]
  PIN rd_out[1559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.785 0.070 722.855 ;
    END
  END rd_out[1559]
  PIN rd_out[1560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 722.925 0.070 722.995 ;
    END
  END rd_out[1560]
  PIN rd_out[1561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.065 0.070 723.135 ;
    END
  END rd_out[1561]
  PIN rd_out[1562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.205 0.070 723.275 ;
    END
  END rd_out[1562]
  PIN rd_out[1563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.345 0.070 723.415 ;
    END
  END rd_out[1563]
  PIN rd_out[1564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.485 0.070 723.555 ;
    END
  END rd_out[1564]
  PIN rd_out[1565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.625 0.070 723.695 ;
    END
  END rd_out[1565]
  PIN rd_out[1566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.765 0.070 723.835 ;
    END
  END rd_out[1566]
  PIN rd_out[1567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 723.905 0.070 723.975 ;
    END
  END rd_out[1567]
  PIN rd_out[1568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.045 0.070 724.115 ;
    END
  END rd_out[1568]
  PIN rd_out[1569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.185 0.070 724.255 ;
    END
  END rd_out[1569]
  PIN rd_out[1570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.325 0.070 724.395 ;
    END
  END rd_out[1570]
  PIN rd_out[1571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.465 0.070 724.535 ;
    END
  END rd_out[1571]
  PIN rd_out[1572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.605 0.070 724.675 ;
    END
  END rd_out[1572]
  PIN rd_out[1573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.745 0.070 724.815 ;
    END
  END rd_out[1573]
  PIN rd_out[1574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 724.885 0.070 724.955 ;
    END
  END rd_out[1574]
  PIN rd_out[1575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.025 0.070 725.095 ;
    END
  END rd_out[1575]
  PIN rd_out[1576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.165 0.070 725.235 ;
    END
  END rd_out[1576]
  PIN rd_out[1577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.305 0.070 725.375 ;
    END
  END rd_out[1577]
  PIN rd_out[1578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.445 0.070 725.515 ;
    END
  END rd_out[1578]
  PIN rd_out[1579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.585 0.070 725.655 ;
    END
  END rd_out[1579]
  PIN rd_out[1580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.725 0.070 725.795 ;
    END
  END rd_out[1580]
  PIN rd_out[1581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 725.865 0.070 725.935 ;
    END
  END rd_out[1581]
  PIN rd_out[1582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.005 0.070 726.075 ;
    END
  END rd_out[1582]
  PIN rd_out[1583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.145 0.070 726.215 ;
    END
  END rd_out[1583]
  PIN rd_out[1584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.285 0.070 726.355 ;
    END
  END rd_out[1584]
  PIN rd_out[1585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.425 0.070 726.495 ;
    END
  END rd_out[1585]
  PIN rd_out[1586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.565 0.070 726.635 ;
    END
  END rd_out[1586]
  PIN rd_out[1587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.705 0.070 726.775 ;
    END
  END rd_out[1587]
  PIN rd_out[1588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.845 0.070 726.915 ;
    END
  END rd_out[1588]
  PIN rd_out[1589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 726.985 0.070 727.055 ;
    END
  END rd_out[1589]
  PIN rd_out[1590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.125 0.070 727.195 ;
    END
  END rd_out[1590]
  PIN rd_out[1591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.265 0.070 727.335 ;
    END
  END rd_out[1591]
  PIN rd_out[1592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.405 0.070 727.475 ;
    END
  END rd_out[1592]
  PIN rd_out[1593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.545 0.070 727.615 ;
    END
  END rd_out[1593]
  PIN rd_out[1594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.685 0.070 727.755 ;
    END
  END rd_out[1594]
  PIN rd_out[1595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.825 0.070 727.895 ;
    END
  END rd_out[1595]
  PIN rd_out[1596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 727.965 0.070 728.035 ;
    END
  END rd_out[1596]
  PIN rd_out[1597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.105 0.070 728.175 ;
    END
  END rd_out[1597]
  PIN rd_out[1598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.245 0.070 728.315 ;
    END
  END rd_out[1598]
  PIN rd_out[1599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.385 0.070 728.455 ;
    END
  END rd_out[1599]
  PIN rd_out[1600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.525 0.070 728.595 ;
    END
  END rd_out[1600]
  PIN rd_out[1601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.665 0.070 728.735 ;
    END
  END rd_out[1601]
  PIN rd_out[1602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.805 0.070 728.875 ;
    END
  END rd_out[1602]
  PIN rd_out[1603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 728.945 0.070 729.015 ;
    END
  END rd_out[1603]
  PIN rd_out[1604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.085 0.070 729.155 ;
    END
  END rd_out[1604]
  PIN rd_out[1605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.225 0.070 729.295 ;
    END
  END rd_out[1605]
  PIN rd_out[1606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.365 0.070 729.435 ;
    END
  END rd_out[1606]
  PIN rd_out[1607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.505 0.070 729.575 ;
    END
  END rd_out[1607]
  PIN rd_out[1608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.645 0.070 729.715 ;
    END
  END rd_out[1608]
  PIN rd_out[1609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.785 0.070 729.855 ;
    END
  END rd_out[1609]
  PIN rd_out[1610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 729.925 0.070 729.995 ;
    END
  END rd_out[1610]
  PIN rd_out[1611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.065 0.070 730.135 ;
    END
  END rd_out[1611]
  PIN rd_out[1612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.205 0.070 730.275 ;
    END
  END rd_out[1612]
  PIN rd_out[1613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.345 0.070 730.415 ;
    END
  END rd_out[1613]
  PIN rd_out[1614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.485 0.070 730.555 ;
    END
  END rd_out[1614]
  PIN rd_out[1615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.625 0.070 730.695 ;
    END
  END rd_out[1615]
  PIN rd_out[1616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.765 0.070 730.835 ;
    END
  END rd_out[1616]
  PIN rd_out[1617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 730.905 0.070 730.975 ;
    END
  END rd_out[1617]
  PIN rd_out[1618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.045 0.070 731.115 ;
    END
  END rd_out[1618]
  PIN rd_out[1619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.185 0.070 731.255 ;
    END
  END rd_out[1619]
  PIN rd_out[1620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.325 0.070 731.395 ;
    END
  END rd_out[1620]
  PIN rd_out[1621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.465 0.070 731.535 ;
    END
  END rd_out[1621]
  PIN rd_out[1622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.605 0.070 731.675 ;
    END
  END rd_out[1622]
  PIN rd_out[1623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.745 0.070 731.815 ;
    END
  END rd_out[1623]
  PIN rd_out[1624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 731.885 0.070 731.955 ;
    END
  END rd_out[1624]
  PIN rd_out[1625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.025 0.070 732.095 ;
    END
  END rd_out[1625]
  PIN rd_out[1626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.165 0.070 732.235 ;
    END
  END rd_out[1626]
  PIN rd_out[1627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.305 0.070 732.375 ;
    END
  END rd_out[1627]
  PIN rd_out[1628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.445 0.070 732.515 ;
    END
  END rd_out[1628]
  PIN rd_out[1629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.585 0.070 732.655 ;
    END
  END rd_out[1629]
  PIN rd_out[1630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.725 0.070 732.795 ;
    END
  END rd_out[1630]
  PIN rd_out[1631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 732.865 0.070 732.935 ;
    END
  END rd_out[1631]
  PIN rd_out[1632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.005 0.070 733.075 ;
    END
  END rd_out[1632]
  PIN rd_out[1633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.145 0.070 733.215 ;
    END
  END rd_out[1633]
  PIN rd_out[1634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.285 0.070 733.355 ;
    END
  END rd_out[1634]
  PIN rd_out[1635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.425 0.070 733.495 ;
    END
  END rd_out[1635]
  PIN rd_out[1636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.565 0.070 733.635 ;
    END
  END rd_out[1636]
  PIN rd_out[1637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.705 0.070 733.775 ;
    END
  END rd_out[1637]
  PIN rd_out[1638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.845 0.070 733.915 ;
    END
  END rd_out[1638]
  PIN rd_out[1639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 733.985 0.070 734.055 ;
    END
  END rd_out[1639]
  PIN rd_out[1640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.125 0.070 734.195 ;
    END
  END rd_out[1640]
  PIN rd_out[1641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.265 0.070 734.335 ;
    END
  END rd_out[1641]
  PIN rd_out[1642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.405 0.070 734.475 ;
    END
  END rd_out[1642]
  PIN rd_out[1643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.545 0.070 734.615 ;
    END
  END rd_out[1643]
  PIN rd_out[1644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.685 0.070 734.755 ;
    END
  END rd_out[1644]
  PIN rd_out[1645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.825 0.070 734.895 ;
    END
  END rd_out[1645]
  PIN rd_out[1646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 734.965 0.070 735.035 ;
    END
  END rd_out[1646]
  PIN rd_out[1647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.105 0.070 735.175 ;
    END
  END rd_out[1647]
  PIN rd_out[1648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.245 0.070 735.315 ;
    END
  END rd_out[1648]
  PIN rd_out[1649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.385 0.070 735.455 ;
    END
  END rd_out[1649]
  PIN rd_out[1650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.525 0.070 735.595 ;
    END
  END rd_out[1650]
  PIN rd_out[1651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.665 0.070 735.735 ;
    END
  END rd_out[1651]
  PIN rd_out[1652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.805 0.070 735.875 ;
    END
  END rd_out[1652]
  PIN rd_out[1653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 735.945 0.070 736.015 ;
    END
  END rd_out[1653]
  PIN rd_out[1654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.085 0.070 736.155 ;
    END
  END rd_out[1654]
  PIN rd_out[1655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.225 0.070 736.295 ;
    END
  END rd_out[1655]
  PIN rd_out[1656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.365 0.070 736.435 ;
    END
  END rd_out[1656]
  PIN rd_out[1657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.505 0.070 736.575 ;
    END
  END rd_out[1657]
  PIN rd_out[1658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.645 0.070 736.715 ;
    END
  END rd_out[1658]
  PIN rd_out[1659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.785 0.070 736.855 ;
    END
  END rd_out[1659]
  PIN rd_out[1660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 736.925 0.070 736.995 ;
    END
  END rd_out[1660]
  PIN rd_out[1661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.065 0.070 737.135 ;
    END
  END rd_out[1661]
  PIN rd_out[1662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.205 0.070 737.275 ;
    END
  END rd_out[1662]
  PIN rd_out[1663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.345 0.070 737.415 ;
    END
  END rd_out[1663]
  PIN rd_out[1664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.485 0.070 737.555 ;
    END
  END rd_out[1664]
  PIN rd_out[1665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.625 0.070 737.695 ;
    END
  END rd_out[1665]
  PIN rd_out[1666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.765 0.070 737.835 ;
    END
  END rd_out[1666]
  PIN rd_out[1667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 737.905 0.070 737.975 ;
    END
  END rd_out[1667]
  PIN rd_out[1668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.045 0.070 738.115 ;
    END
  END rd_out[1668]
  PIN rd_out[1669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.185 0.070 738.255 ;
    END
  END rd_out[1669]
  PIN rd_out[1670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.325 0.070 738.395 ;
    END
  END rd_out[1670]
  PIN rd_out[1671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.465 0.070 738.535 ;
    END
  END rd_out[1671]
  PIN rd_out[1672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.605 0.070 738.675 ;
    END
  END rd_out[1672]
  PIN rd_out[1673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.745 0.070 738.815 ;
    END
  END rd_out[1673]
  PIN rd_out[1674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 738.885 0.070 738.955 ;
    END
  END rd_out[1674]
  PIN rd_out[1675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.025 0.070 739.095 ;
    END
  END rd_out[1675]
  PIN rd_out[1676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.165 0.070 739.235 ;
    END
  END rd_out[1676]
  PIN rd_out[1677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.305 0.070 739.375 ;
    END
  END rd_out[1677]
  PIN rd_out[1678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.445 0.070 739.515 ;
    END
  END rd_out[1678]
  PIN rd_out[1679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.585 0.070 739.655 ;
    END
  END rd_out[1679]
  PIN rd_out[1680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.725 0.070 739.795 ;
    END
  END rd_out[1680]
  PIN rd_out[1681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 739.865 0.070 739.935 ;
    END
  END rd_out[1681]
  PIN rd_out[1682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.005 0.070 740.075 ;
    END
  END rd_out[1682]
  PIN rd_out[1683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.145 0.070 740.215 ;
    END
  END rd_out[1683]
  PIN rd_out[1684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.285 0.070 740.355 ;
    END
  END rd_out[1684]
  PIN rd_out[1685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.425 0.070 740.495 ;
    END
  END rd_out[1685]
  PIN rd_out[1686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.565 0.070 740.635 ;
    END
  END rd_out[1686]
  PIN rd_out[1687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.705 0.070 740.775 ;
    END
  END rd_out[1687]
  PIN rd_out[1688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.845 0.070 740.915 ;
    END
  END rd_out[1688]
  PIN rd_out[1689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 740.985 0.070 741.055 ;
    END
  END rd_out[1689]
  PIN rd_out[1690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.125 0.070 741.195 ;
    END
  END rd_out[1690]
  PIN rd_out[1691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.265 0.070 741.335 ;
    END
  END rd_out[1691]
  PIN rd_out[1692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.405 0.070 741.475 ;
    END
  END rd_out[1692]
  PIN rd_out[1693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.545 0.070 741.615 ;
    END
  END rd_out[1693]
  PIN rd_out[1694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.685 0.070 741.755 ;
    END
  END rd_out[1694]
  PIN rd_out[1695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.825 0.070 741.895 ;
    END
  END rd_out[1695]
  PIN rd_out[1696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 741.965 0.070 742.035 ;
    END
  END rd_out[1696]
  PIN rd_out[1697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.105 0.070 742.175 ;
    END
  END rd_out[1697]
  PIN rd_out[1698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.245 0.070 742.315 ;
    END
  END rd_out[1698]
  PIN rd_out[1699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.385 0.070 742.455 ;
    END
  END rd_out[1699]
  PIN rd_out[1700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.525 0.070 742.595 ;
    END
  END rd_out[1700]
  PIN rd_out[1701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.665 0.070 742.735 ;
    END
  END rd_out[1701]
  PIN rd_out[1702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.805 0.070 742.875 ;
    END
  END rd_out[1702]
  PIN rd_out[1703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 742.945 0.070 743.015 ;
    END
  END rd_out[1703]
  PIN rd_out[1704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.085 0.070 743.155 ;
    END
  END rd_out[1704]
  PIN rd_out[1705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.225 0.070 743.295 ;
    END
  END rd_out[1705]
  PIN rd_out[1706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.365 0.070 743.435 ;
    END
  END rd_out[1706]
  PIN rd_out[1707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.505 0.070 743.575 ;
    END
  END rd_out[1707]
  PIN rd_out[1708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.645 0.070 743.715 ;
    END
  END rd_out[1708]
  PIN rd_out[1709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.785 0.070 743.855 ;
    END
  END rd_out[1709]
  PIN rd_out[1710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 743.925 0.070 743.995 ;
    END
  END rd_out[1710]
  PIN rd_out[1711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.065 0.070 744.135 ;
    END
  END rd_out[1711]
  PIN rd_out[1712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.205 0.070 744.275 ;
    END
  END rd_out[1712]
  PIN rd_out[1713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.345 0.070 744.415 ;
    END
  END rd_out[1713]
  PIN rd_out[1714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.485 0.070 744.555 ;
    END
  END rd_out[1714]
  PIN rd_out[1715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.625 0.070 744.695 ;
    END
  END rd_out[1715]
  PIN rd_out[1716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.765 0.070 744.835 ;
    END
  END rd_out[1716]
  PIN rd_out[1717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 744.905 0.070 744.975 ;
    END
  END rd_out[1717]
  PIN rd_out[1718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.045 0.070 745.115 ;
    END
  END rd_out[1718]
  PIN rd_out[1719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.185 0.070 745.255 ;
    END
  END rd_out[1719]
  PIN rd_out[1720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.325 0.070 745.395 ;
    END
  END rd_out[1720]
  PIN rd_out[1721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.465 0.070 745.535 ;
    END
  END rd_out[1721]
  PIN rd_out[1722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.605 0.070 745.675 ;
    END
  END rd_out[1722]
  PIN rd_out[1723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.745 0.070 745.815 ;
    END
  END rd_out[1723]
  PIN rd_out[1724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 745.885 0.070 745.955 ;
    END
  END rd_out[1724]
  PIN rd_out[1725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.025 0.070 746.095 ;
    END
  END rd_out[1725]
  PIN rd_out[1726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.165 0.070 746.235 ;
    END
  END rd_out[1726]
  PIN rd_out[1727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.305 0.070 746.375 ;
    END
  END rd_out[1727]
  PIN rd_out[1728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.445 0.070 746.515 ;
    END
  END rd_out[1728]
  PIN rd_out[1729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.585 0.070 746.655 ;
    END
  END rd_out[1729]
  PIN rd_out[1730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.725 0.070 746.795 ;
    END
  END rd_out[1730]
  PIN rd_out[1731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 746.865 0.070 746.935 ;
    END
  END rd_out[1731]
  PIN rd_out[1732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.005 0.070 747.075 ;
    END
  END rd_out[1732]
  PIN rd_out[1733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.145 0.070 747.215 ;
    END
  END rd_out[1733]
  PIN rd_out[1734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.285 0.070 747.355 ;
    END
  END rd_out[1734]
  PIN rd_out[1735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.425 0.070 747.495 ;
    END
  END rd_out[1735]
  PIN rd_out[1736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.565 0.070 747.635 ;
    END
  END rd_out[1736]
  PIN rd_out[1737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.705 0.070 747.775 ;
    END
  END rd_out[1737]
  PIN rd_out[1738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.845 0.070 747.915 ;
    END
  END rd_out[1738]
  PIN rd_out[1739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 747.985 0.070 748.055 ;
    END
  END rd_out[1739]
  PIN rd_out[1740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.125 0.070 748.195 ;
    END
  END rd_out[1740]
  PIN rd_out[1741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.265 0.070 748.335 ;
    END
  END rd_out[1741]
  PIN rd_out[1742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.405 0.070 748.475 ;
    END
  END rd_out[1742]
  PIN rd_out[1743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.545 0.070 748.615 ;
    END
  END rd_out[1743]
  PIN rd_out[1744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.685 0.070 748.755 ;
    END
  END rd_out[1744]
  PIN rd_out[1745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.825 0.070 748.895 ;
    END
  END rd_out[1745]
  PIN rd_out[1746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 748.965 0.070 749.035 ;
    END
  END rd_out[1746]
  PIN rd_out[1747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.105 0.070 749.175 ;
    END
  END rd_out[1747]
  PIN rd_out[1748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.245 0.070 749.315 ;
    END
  END rd_out[1748]
  PIN rd_out[1749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.385 0.070 749.455 ;
    END
  END rd_out[1749]
  PIN rd_out[1750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.525 0.070 749.595 ;
    END
  END rd_out[1750]
  PIN rd_out[1751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.665 0.070 749.735 ;
    END
  END rd_out[1751]
  PIN rd_out[1752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.805 0.070 749.875 ;
    END
  END rd_out[1752]
  PIN rd_out[1753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 749.945 0.070 750.015 ;
    END
  END rd_out[1753]
  PIN rd_out[1754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.085 0.070 750.155 ;
    END
  END rd_out[1754]
  PIN rd_out[1755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.225 0.070 750.295 ;
    END
  END rd_out[1755]
  PIN rd_out[1756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.365 0.070 750.435 ;
    END
  END rd_out[1756]
  PIN rd_out[1757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.505 0.070 750.575 ;
    END
  END rd_out[1757]
  PIN rd_out[1758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.645 0.070 750.715 ;
    END
  END rd_out[1758]
  PIN rd_out[1759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.785 0.070 750.855 ;
    END
  END rd_out[1759]
  PIN rd_out[1760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 750.925 0.070 750.995 ;
    END
  END rd_out[1760]
  PIN rd_out[1761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.065 0.070 751.135 ;
    END
  END rd_out[1761]
  PIN rd_out[1762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.205 0.070 751.275 ;
    END
  END rd_out[1762]
  PIN rd_out[1763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.345 0.070 751.415 ;
    END
  END rd_out[1763]
  PIN rd_out[1764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.485 0.070 751.555 ;
    END
  END rd_out[1764]
  PIN rd_out[1765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.625 0.070 751.695 ;
    END
  END rd_out[1765]
  PIN rd_out[1766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.765 0.070 751.835 ;
    END
  END rd_out[1766]
  PIN rd_out[1767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 751.905 0.070 751.975 ;
    END
  END rd_out[1767]
  PIN rd_out[1768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.045 0.070 752.115 ;
    END
  END rd_out[1768]
  PIN rd_out[1769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.185 0.070 752.255 ;
    END
  END rd_out[1769]
  PIN rd_out[1770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.325 0.070 752.395 ;
    END
  END rd_out[1770]
  PIN rd_out[1771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.465 0.070 752.535 ;
    END
  END rd_out[1771]
  PIN rd_out[1772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.605 0.070 752.675 ;
    END
  END rd_out[1772]
  PIN rd_out[1773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.745 0.070 752.815 ;
    END
  END rd_out[1773]
  PIN rd_out[1774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 752.885 0.070 752.955 ;
    END
  END rd_out[1774]
  PIN rd_out[1775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.025 0.070 753.095 ;
    END
  END rd_out[1775]
  PIN rd_out[1776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.165 0.070 753.235 ;
    END
  END rd_out[1776]
  PIN rd_out[1777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.305 0.070 753.375 ;
    END
  END rd_out[1777]
  PIN rd_out[1778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.445 0.070 753.515 ;
    END
  END rd_out[1778]
  PIN rd_out[1779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.585 0.070 753.655 ;
    END
  END rd_out[1779]
  PIN rd_out[1780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.725 0.070 753.795 ;
    END
  END rd_out[1780]
  PIN rd_out[1781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 753.865 0.070 753.935 ;
    END
  END rd_out[1781]
  PIN rd_out[1782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.005 0.070 754.075 ;
    END
  END rd_out[1782]
  PIN rd_out[1783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.145 0.070 754.215 ;
    END
  END rd_out[1783]
  PIN rd_out[1784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.285 0.070 754.355 ;
    END
  END rd_out[1784]
  PIN rd_out[1785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.425 0.070 754.495 ;
    END
  END rd_out[1785]
  PIN rd_out[1786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.565 0.070 754.635 ;
    END
  END rd_out[1786]
  PIN rd_out[1787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.705 0.070 754.775 ;
    END
  END rd_out[1787]
  PIN rd_out[1788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.845 0.070 754.915 ;
    END
  END rd_out[1788]
  PIN rd_out[1789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 754.985 0.070 755.055 ;
    END
  END rd_out[1789]
  PIN rd_out[1790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.125 0.070 755.195 ;
    END
  END rd_out[1790]
  PIN rd_out[1791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.265 0.070 755.335 ;
    END
  END rd_out[1791]
  PIN rd_out[1792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.405 0.070 755.475 ;
    END
  END rd_out[1792]
  PIN rd_out[1793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.545 0.070 755.615 ;
    END
  END rd_out[1793]
  PIN rd_out[1794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.685 0.070 755.755 ;
    END
  END rd_out[1794]
  PIN rd_out[1795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.825 0.070 755.895 ;
    END
  END rd_out[1795]
  PIN rd_out[1796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 755.965 0.070 756.035 ;
    END
  END rd_out[1796]
  PIN rd_out[1797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.105 0.070 756.175 ;
    END
  END rd_out[1797]
  PIN rd_out[1798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.245 0.070 756.315 ;
    END
  END rd_out[1798]
  PIN rd_out[1799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.385 0.070 756.455 ;
    END
  END rd_out[1799]
  PIN rd_out[1800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.525 0.070 756.595 ;
    END
  END rd_out[1800]
  PIN rd_out[1801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.665 0.070 756.735 ;
    END
  END rd_out[1801]
  PIN rd_out[1802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.805 0.070 756.875 ;
    END
  END rd_out[1802]
  PIN rd_out[1803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 756.945 0.070 757.015 ;
    END
  END rd_out[1803]
  PIN rd_out[1804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.085 0.070 757.155 ;
    END
  END rd_out[1804]
  PIN rd_out[1805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.225 0.070 757.295 ;
    END
  END rd_out[1805]
  PIN rd_out[1806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.365 0.070 757.435 ;
    END
  END rd_out[1806]
  PIN rd_out[1807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.505 0.070 757.575 ;
    END
  END rd_out[1807]
  PIN rd_out[1808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.645 0.070 757.715 ;
    END
  END rd_out[1808]
  PIN rd_out[1809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.785 0.070 757.855 ;
    END
  END rd_out[1809]
  PIN rd_out[1810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 757.925 0.070 757.995 ;
    END
  END rd_out[1810]
  PIN rd_out[1811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.065 0.070 758.135 ;
    END
  END rd_out[1811]
  PIN rd_out[1812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.205 0.070 758.275 ;
    END
  END rd_out[1812]
  PIN rd_out[1813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.345 0.070 758.415 ;
    END
  END rd_out[1813]
  PIN rd_out[1814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.485 0.070 758.555 ;
    END
  END rd_out[1814]
  PIN rd_out[1815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.625 0.070 758.695 ;
    END
  END rd_out[1815]
  PIN rd_out[1816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.765 0.070 758.835 ;
    END
  END rd_out[1816]
  PIN rd_out[1817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 758.905 0.070 758.975 ;
    END
  END rd_out[1817]
  PIN rd_out[1818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.045 0.070 759.115 ;
    END
  END rd_out[1818]
  PIN rd_out[1819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.185 0.070 759.255 ;
    END
  END rd_out[1819]
  PIN rd_out[1820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.325 0.070 759.395 ;
    END
  END rd_out[1820]
  PIN rd_out[1821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.465 0.070 759.535 ;
    END
  END rd_out[1821]
  PIN rd_out[1822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.605 0.070 759.675 ;
    END
  END rd_out[1822]
  PIN rd_out[1823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.745 0.070 759.815 ;
    END
  END rd_out[1823]
  PIN rd_out[1824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 759.885 0.070 759.955 ;
    END
  END rd_out[1824]
  PIN rd_out[1825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.025 0.070 760.095 ;
    END
  END rd_out[1825]
  PIN rd_out[1826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.165 0.070 760.235 ;
    END
  END rd_out[1826]
  PIN rd_out[1827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.305 0.070 760.375 ;
    END
  END rd_out[1827]
  PIN rd_out[1828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.445 0.070 760.515 ;
    END
  END rd_out[1828]
  PIN rd_out[1829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.585 0.070 760.655 ;
    END
  END rd_out[1829]
  PIN rd_out[1830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.725 0.070 760.795 ;
    END
  END rd_out[1830]
  PIN rd_out[1831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 760.865 0.070 760.935 ;
    END
  END rd_out[1831]
  PIN rd_out[1832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.005 0.070 761.075 ;
    END
  END rd_out[1832]
  PIN rd_out[1833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.145 0.070 761.215 ;
    END
  END rd_out[1833]
  PIN rd_out[1834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.285 0.070 761.355 ;
    END
  END rd_out[1834]
  PIN rd_out[1835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.425 0.070 761.495 ;
    END
  END rd_out[1835]
  PIN rd_out[1836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.565 0.070 761.635 ;
    END
  END rd_out[1836]
  PIN rd_out[1837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.705 0.070 761.775 ;
    END
  END rd_out[1837]
  PIN rd_out[1838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.845 0.070 761.915 ;
    END
  END rd_out[1838]
  PIN rd_out[1839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 761.985 0.070 762.055 ;
    END
  END rd_out[1839]
  PIN rd_out[1840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.125 0.070 762.195 ;
    END
  END rd_out[1840]
  PIN rd_out[1841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.265 0.070 762.335 ;
    END
  END rd_out[1841]
  PIN rd_out[1842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.405 0.070 762.475 ;
    END
  END rd_out[1842]
  PIN rd_out[1843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.545 0.070 762.615 ;
    END
  END rd_out[1843]
  PIN rd_out[1844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.685 0.070 762.755 ;
    END
  END rd_out[1844]
  PIN rd_out[1845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.825 0.070 762.895 ;
    END
  END rd_out[1845]
  PIN rd_out[1846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 762.965 0.070 763.035 ;
    END
  END rd_out[1846]
  PIN rd_out[1847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.105 0.070 763.175 ;
    END
  END rd_out[1847]
  PIN rd_out[1848]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.245 0.070 763.315 ;
    END
  END rd_out[1848]
  PIN rd_out[1849]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.385 0.070 763.455 ;
    END
  END rd_out[1849]
  PIN rd_out[1850]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.525 0.070 763.595 ;
    END
  END rd_out[1850]
  PIN rd_out[1851]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.665 0.070 763.735 ;
    END
  END rd_out[1851]
  PIN rd_out[1852]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.805 0.070 763.875 ;
    END
  END rd_out[1852]
  PIN rd_out[1853]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 763.945 0.070 764.015 ;
    END
  END rd_out[1853]
  PIN rd_out[1854]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.085 0.070 764.155 ;
    END
  END rd_out[1854]
  PIN rd_out[1855]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.225 0.070 764.295 ;
    END
  END rd_out[1855]
  PIN rd_out[1856]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.365 0.070 764.435 ;
    END
  END rd_out[1856]
  PIN rd_out[1857]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.505 0.070 764.575 ;
    END
  END rd_out[1857]
  PIN rd_out[1858]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.645 0.070 764.715 ;
    END
  END rd_out[1858]
  PIN rd_out[1859]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.785 0.070 764.855 ;
    END
  END rd_out[1859]
  PIN rd_out[1860]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 764.925 0.070 764.995 ;
    END
  END rd_out[1860]
  PIN rd_out[1861]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.065 0.070 765.135 ;
    END
  END rd_out[1861]
  PIN rd_out[1862]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.205 0.070 765.275 ;
    END
  END rd_out[1862]
  PIN rd_out[1863]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.345 0.070 765.415 ;
    END
  END rd_out[1863]
  PIN rd_out[1864]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.485 0.070 765.555 ;
    END
  END rd_out[1864]
  PIN rd_out[1865]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.625 0.070 765.695 ;
    END
  END rd_out[1865]
  PIN rd_out[1866]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.765 0.070 765.835 ;
    END
  END rd_out[1866]
  PIN rd_out[1867]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 765.905 0.070 765.975 ;
    END
  END rd_out[1867]
  PIN rd_out[1868]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.045 0.070 766.115 ;
    END
  END rd_out[1868]
  PIN rd_out[1869]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.185 0.070 766.255 ;
    END
  END rd_out[1869]
  PIN rd_out[1870]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.325 0.070 766.395 ;
    END
  END rd_out[1870]
  PIN rd_out[1871]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.465 0.070 766.535 ;
    END
  END rd_out[1871]
  PIN rd_out[1872]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.605 0.070 766.675 ;
    END
  END rd_out[1872]
  PIN rd_out[1873]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.745 0.070 766.815 ;
    END
  END rd_out[1873]
  PIN rd_out[1874]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 766.885 0.070 766.955 ;
    END
  END rd_out[1874]
  PIN rd_out[1875]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.025 0.070 767.095 ;
    END
  END rd_out[1875]
  PIN rd_out[1876]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.165 0.070 767.235 ;
    END
  END rd_out[1876]
  PIN rd_out[1877]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.305 0.070 767.375 ;
    END
  END rd_out[1877]
  PIN rd_out[1878]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.445 0.070 767.515 ;
    END
  END rd_out[1878]
  PIN rd_out[1879]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.585 0.070 767.655 ;
    END
  END rd_out[1879]
  PIN rd_out[1880]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.725 0.070 767.795 ;
    END
  END rd_out[1880]
  PIN rd_out[1881]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 767.865 0.070 767.935 ;
    END
  END rd_out[1881]
  PIN rd_out[1882]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.005 0.070 768.075 ;
    END
  END rd_out[1882]
  PIN rd_out[1883]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.145 0.070 768.215 ;
    END
  END rd_out[1883]
  PIN rd_out[1884]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.285 0.070 768.355 ;
    END
  END rd_out[1884]
  PIN rd_out[1885]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.425 0.070 768.495 ;
    END
  END rd_out[1885]
  PIN rd_out[1886]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.565 0.070 768.635 ;
    END
  END rd_out[1886]
  PIN rd_out[1887]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.705 0.070 768.775 ;
    END
  END rd_out[1887]
  PIN rd_out[1888]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.845 0.070 768.915 ;
    END
  END rd_out[1888]
  PIN rd_out[1889]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 768.985 0.070 769.055 ;
    END
  END rd_out[1889]
  PIN rd_out[1890]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.125 0.070 769.195 ;
    END
  END rd_out[1890]
  PIN rd_out[1891]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.265 0.070 769.335 ;
    END
  END rd_out[1891]
  PIN rd_out[1892]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.405 0.070 769.475 ;
    END
  END rd_out[1892]
  PIN rd_out[1893]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.545 0.070 769.615 ;
    END
  END rd_out[1893]
  PIN rd_out[1894]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.685 0.070 769.755 ;
    END
  END rd_out[1894]
  PIN rd_out[1895]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.825 0.070 769.895 ;
    END
  END rd_out[1895]
  PIN rd_out[1896]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 769.965 0.070 770.035 ;
    END
  END rd_out[1896]
  PIN rd_out[1897]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.105 0.070 770.175 ;
    END
  END rd_out[1897]
  PIN rd_out[1898]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.245 0.070 770.315 ;
    END
  END rd_out[1898]
  PIN rd_out[1899]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.385 0.070 770.455 ;
    END
  END rd_out[1899]
  PIN rd_out[1900]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.525 0.070 770.595 ;
    END
  END rd_out[1900]
  PIN rd_out[1901]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.665 0.070 770.735 ;
    END
  END rd_out[1901]
  PIN rd_out[1902]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.805 0.070 770.875 ;
    END
  END rd_out[1902]
  PIN rd_out[1903]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 770.945 0.070 771.015 ;
    END
  END rd_out[1903]
  PIN rd_out[1904]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.085 0.070 771.155 ;
    END
  END rd_out[1904]
  PIN rd_out[1905]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.225 0.070 771.295 ;
    END
  END rd_out[1905]
  PIN rd_out[1906]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.365 0.070 771.435 ;
    END
  END rd_out[1906]
  PIN rd_out[1907]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.505 0.070 771.575 ;
    END
  END rd_out[1907]
  PIN rd_out[1908]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.645 0.070 771.715 ;
    END
  END rd_out[1908]
  PIN rd_out[1909]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.785 0.070 771.855 ;
    END
  END rd_out[1909]
  PIN rd_out[1910]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 771.925 0.070 771.995 ;
    END
  END rd_out[1910]
  PIN rd_out[1911]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.065 0.070 772.135 ;
    END
  END rd_out[1911]
  PIN rd_out[1912]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.205 0.070 772.275 ;
    END
  END rd_out[1912]
  PIN rd_out[1913]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.345 0.070 772.415 ;
    END
  END rd_out[1913]
  PIN rd_out[1914]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.485 0.070 772.555 ;
    END
  END rd_out[1914]
  PIN rd_out[1915]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.625 0.070 772.695 ;
    END
  END rd_out[1915]
  PIN rd_out[1916]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.765 0.070 772.835 ;
    END
  END rd_out[1916]
  PIN rd_out[1917]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 772.905 0.070 772.975 ;
    END
  END rd_out[1917]
  PIN rd_out[1918]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.045 0.070 773.115 ;
    END
  END rd_out[1918]
  PIN rd_out[1919]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.185 0.070 773.255 ;
    END
  END rd_out[1919]
  PIN rd_out[1920]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.325 0.070 773.395 ;
    END
  END rd_out[1920]
  PIN rd_out[1921]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.465 0.070 773.535 ;
    END
  END rd_out[1921]
  PIN rd_out[1922]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.605 0.070 773.675 ;
    END
  END rd_out[1922]
  PIN rd_out[1923]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.745 0.070 773.815 ;
    END
  END rd_out[1923]
  PIN rd_out[1924]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 773.885 0.070 773.955 ;
    END
  END rd_out[1924]
  PIN rd_out[1925]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 774.025 0.070 774.095 ;
    END
  END rd_out[1925]
  PIN rd_out[1926]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 774.165 0.070 774.235 ;
    END
  END rd_out[1926]
  PIN rd_out[1927]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 774.305 0.070 774.375 ;
    END
  END rd_out[1927]
  PIN rd_out[1928]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 774.445 0.070 774.515 ;
    END
  END rd_out[1928]
  PIN rd_out[1929]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 774.585 0.070 774.655 ;
    END
  END rd_out[1929]
  PIN rd_out[1930]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 774.725 0.070 774.795 ;
    END
  END rd_out[1930]
  PIN rd_out[1931]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 774.865 0.070 774.935 ;
    END
  END rd_out[1931]
  PIN rd_out[1932]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.005 0.070 775.075 ;
    END
  END rd_out[1932]
  PIN rd_out[1933]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.145 0.070 775.215 ;
    END
  END rd_out[1933]
  PIN rd_out[1934]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.285 0.070 775.355 ;
    END
  END rd_out[1934]
  PIN rd_out[1935]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.425 0.070 775.495 ;
    END
  END rd_out[1935]
  PIN rd_out[1936]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.565 0.070 775.635 ;
    END
  END rd_out[1936]
  PIN rd_out[1937]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.705 0.070 775.775 ;
    END
  END rd_out[1937]
  PIN rd_out[1938]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.845 0.070 775.915 ;
    END
  END rd_out[1938]
  PIN rd_out[1939]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 775.985 0.070 776.055 ;
    END
  END rd_out[1939]
  PIN rd_out[1940]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.125 0.070 776.195 ;
    END
  END rd_out[1940]
  PIN rd_out[1941]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.265 0.070 776.335 ;
    END
  END rd_out[1941]
  PIN rd_out[1942]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.405 0.070 776.475 ;
    END
  END rd_out[1942]
  PIN rd_out[1943]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.545 0.070 776.615 ;
    END
  END rd_out[1943]
  PIN rd_out[1944]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.685 0.070 776.755 ;
    END
  END rd_out[1944]
  PIN rd_out[1945]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.825 0.070 776.895 ;
    END
  END rd_out[1945]
  PIN rd_out[1946]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 776.965 0.070 777.035 ;
    END
  END rd_out[1946]
  PIN rd_out[1947]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.105 0.070 777.175 ;
    END
  END rd_out[1947]
  PIN rd_out[1948]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.245 0.070 777.315 ;
    END
  END rd_out[1948]
  PIN rd_out[1949]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.385 0.070 777.455 ;
    END
  END rd_out[1949]
  PIN rd_out[1950]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.525 0.070 777.595 ;
    END
  END rd_out[1950]
  PIN rd_out[1951]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.665 0.070 777.735 ;
    END
  END rd_out[1951]
  PIN rd_out[1952]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.805 0.070 777.875 ;
    END
  END rd_out[1952]
  PIN rd_out[1953]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 777.945 0.070 778.015 ;
    END
  END rd_out[1953]
  PIN rd_out[1954]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.085 0.070 778.155 ;
    END
  END rd_out[1954]
  PIN rd_out[1955]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.225 0.070 778.295 ;
    END
  END rd_out[1955]
  PIN rd_out[1956]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.365 0.070 778.435 ;
    END
  END rd_out[1956]
  PIN rd_out[1957]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.505 0.070 778.575 ;
    END
  END rd_out[1957]
  PIN rd_out[1958]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.645 0.070 778.715 ;
    END
  END rd_out[1958]
  PIN rd_out[1959]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.785 0.070 778.855 ;
    END
  END rd_out[1959]
  PIN rd_out[1960]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 778.925 0.070 778.995 ;
    END
  END rd_out[1960]
  PIN rd_out[1961]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 779.065 0.070 779.135 ;
    END
  END rd_out[1961]
  PIN rd_out[1962]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 779.205 0.070 779.275 ;
    END
  END rd_out[1962]
  PIN rd_out[1963]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 779.345 0.070 779.415 ;
    END
  END rd_out[1963]
  PIN rd_out[1964]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 779.485 0.070 779.555 ;
    END
  END rd_out[1964]
  PIN rd_out[1965]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 779.625 0.070 779.695 ;
    END
  END rd_out[1965]
  PIN rd_out[1966]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 779.765 0.070 779.835 ;
    END
  END rd_out[1966]
  PIN rd_out[1967]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 779.905 0.070 779.975 ;
    END
  END rd_out[1967]
  PIN rd_out[1968]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.045 0.070 780.115 ;
    END
  END rd_out[1968]
  PIN rd_out[1969]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.185 0.070 780.255 ;
    END
  END rd_out[1969]
  PIN rd_out[1970]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.325 0.070 780.395 ;
    END
  END rd_out[1970]
  PIN rd_out[1971]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.465 0.070 780.535 ;
    END
  END rd_out[1971]
  PIN rd_out[1972]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.605 0.070 780.675 ;
    END
  END rd_out[1972]
  PIN rd_out[1973]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.745 0.070 780.815 ;
    END
  END rd_out[1973]
  PIN rd_out[1974]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 780.885 0.070 780.955 ;
    END
  END rd_out[1974]
  PIN rd_out[1975]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.025 0.070 781.095 ;
    END
  END rd_out[1975]
  PIN rd_out[1976]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.165 0.070 781.235 ;
    END
  END rd_out[1976]
  PIN rd_out[1977]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.305 0.070 781.375 ;
    END
  END rd_out[1977]
  PIN rd_out[1978]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.445 0.070 781.515 ;
    END
  END rd_out[1978]
  PIN rd_out[1979]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.585 0.070 781.655 ;
    END
  END rd_out[1979]
  PIN rd_out[1980]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.725 0.070 781.795 ;
    END
  END rd_out[1980]
  PIN rd_out[1981]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 781.865 0.070 781.935 ;
    END
  END rd_out[1981]
  PIN rd_out[1982]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.005 0.070 782.075 ;
    END
  END rd_out[1982]
  PIN rd_out[1983]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.145 0.070 782.215 ;
    END
  END rd_out[1983]
  PIN rd_out[1984]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.285 0.070 782.355 ;
    END
  END rd_out[1984]
  PIN rd_out[1985]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.425 0.070 782.495 ;
    END
  END rd_out[1985]
  PIN rd_out[1986]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.565 0.070 782.635 ;
    END
  END rd_out[1986]
  PIN rd_out[1987]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.705 0.070 782.775 ;
    END
  END rd_out[1987]
  PIN rd_out[1988]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.845 0.070 782.915 ;
    END
  END rd_out[1988]
  PIN rd_out[1989]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 782.985 0.070 783.055 ;
    END
  END rd_out[1989]
  PIN rd_out[1990]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.125 0.070 783.195 ;
    END
  END rd_out[1990]
  PIN rd_out[1991]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.265 0.070 783.335 ;
    END
  END rd_out[1991]
  PIN rd_out[1992]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.405 0.070 783.475 ;
    END
  END rd_out[1992]
  PIN rd_out[1993]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.545 0.070 783.615 ;
    END
  END rd_out[1993]
  PIN rd_out[1994]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.685 0.070 783.755 ;
    END
  END rd_out[1994]
  PIN rd_out[1995]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.825 0.070 783.895 ;
    END
  END rd_out[1995]
  PIN rd_out[1996]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 783.965 0.070 784.035 ;
    END
  END rd_out[1996]
  PIN rd_out[1997]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 784.105 0.070 784.175 ;
    END
  END rd_out[1997]
  PIN rd_out[1998]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 784.245 0.070 784.315 ;
    END
  END rd_out[1998]
  PIN rd_out[1999]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 784.385 0.070 784.455 ;
    END
  END rd_out[1999]
  PIN rd_out[2000]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 784.525 0.070 784.595 ;
    END
  END rd_out[2000]
  PIN rd_out[2001]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 784.665 0.070 784.735 ;
    END
  END rd_out[2001]
  PIN rd_out[2002]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 784.805 0.070 784.875 ;
    END
  END rd_out[2002]
  PIN rd_out[2003]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 784.945 0.070 785.015 ;
    END
  END rd_out[2003]
  PIN rd_out[2004]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.085 0.070 785.155 ;
    END
  END rd_out[2004]
  PIN rd_out[2005]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.225 0.070 785.295 ;
    END
  END rd_out[2005]
  PIN rd_out[2006]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.365 0.070 785.435 ;
    END
  END rd_out[2006]
  PIN rd_out[2007]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.505 0.070 785.575 ;
    END
  END rd_out[2007]
  PIN rd_out[2008]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.645 0.070 785.715 ;
    END
  END rd_out[2008]
  PIN rd_out[2009]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.785 0.070 785.855 ;
    END
  END rd_out[2009]
  PIN rd_out[2010]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 785.925 0.070 785.995 ;
    END
  END rd_out[2010]
  PIN rd_out[2011]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.065 0.070 786.135 ;
    END
  END rd_out[2011]
  PIN rd_out[2012]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.205 0.070 786.275 ;
    END
  END rd_out[2012]
  PIN rd_out[2013]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.345 0.070 786.415 ;
    END
  END rd_out[2013]
  PIN rd_out[2014]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.485 0.070 786.555 ;
    END
  END rd_out[2014]
  PIN rd_out[2015]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.625 0.070 786.695 ;
    END
  END rd_out[2015]
  PIN rd_out[2016]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.765 0.070 786.835 ;
    END
  END rd_out[2016]
  PIN rd_out[2017]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 786.905 0.070 786.975 ;
    END
  END rd_out[2017]
  PIN rd_out[2018]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.045 0.070 787.115 ;
    END
  END rd_out[2018]
  PIN rd_out[2019]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.185 0.070 787.255 ;
    END
  END rd_out[2019]
  PIN rd_out[2020]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.325 0.070 787.395 ;
    END
  END rd_out[2020]
  PIN rd_out[2021]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.465 0.070 787.535 ;
    END
  END rd_out[2021]
  PIN rd_out[2022]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.605 0.070 787.675 ;
    END
  END rd_out[2022]
  PIN rd_out[2023]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.745 0.070 787.815 ;
    END
  END rd_out[2023]
  PIN rd_out[2024]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 787.885 0.070 787.955 ;
    END
  END rd_out[2024]
  PIN rd_out[2025]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 788.025 0.070 788.095 ;
    END
  END rd_out[2025]
  PIN rd_out[2026]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 788.165 0.070 788.235 ;
    END
  END rd_out[2026]
  PIN rd_out[2027]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 788.305 0.070 788.375 ;
    END
  END rd_out[2027]
  PIN rd_out[2028]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 788.445 0.070 788.515 ;
    END
  END rd_out[2028]
  PIN rd_out[2029]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 788.585 0.070 788.655 ;
    END
  END rd_out[2029]
  PIN rd_out[2030]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 788.725 0.070 788.795 ;
    END
  END rd_out[2030]
  PIN rd_out[2031]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 788.865 0.070 788.935 ;
    END
  END rd_out[2031]
  PIN rd_out[2032]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.005 0.070 789.075 ;
    END
  END rd_out[2032]
  PIN rd_out[2033]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.145 0.070 789.215 ;
    END
  END rd_out[2033]
  PIN rd_out[2034]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.285 0.070 789.355 ;
    END
  END rd_out[2034]
  PIN rd_out[2035]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.425 0.070 789.495 ;
    END
  END rd_out[2035]
  PIN rd_out[2036]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.565 0.070 789.635 ;
    END
  END rd_out[2036]
  PIN rd_out[2037]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.705 0.070 789.775 ;
    END
  END rd_out[2037]
  PIN rd_out[2038]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.845 0.070 789.915 ;
    END
  END rd_out[2038]
  PIN rd_out[2039]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 789.985 0.070 790.055 ;
    END
  END rd_out[2039]
  PIN rd_out[2040]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.125 0.070 790.195 ;
    END
  END rd_out[2040]
  PIN rd_out[2041]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.265 0.070 790.335 ;
    END
  END rd_out[2041]
  PIN rd_out[2042]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.405 0.070 790.475 ;
    END
  END rd_out[2042]
  PIN rd_out[2043]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.545 0.070 790.615 ;
    END
  END rd_out[2043]
  PIN rd_out[2044]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.685 0.070 790.755 ;
    END
  END rd_out[2044]
  PIN rd_out[2045]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.825 0.070 790.895 ;
    END
  END rd_out[2045]
  PIN rd_out[2046]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 790.965 0.070 791.035 ;
    END
  END rd_out[2046]
  PIN rd_out[2047]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.105 0.070 791.175 ;
    END
  END rd_out[2047]
  PIN rd_out[2048]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.245 0.070 791.315 ;
    END
  END rd_out[2048]
  PIN rd_out[2049]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.385 0.070 791.455 ;
    END
  END rd_out[2049]
  PIN rd_out[2050]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.525 0.070 791.595 ;
    END
  END rd_out[2050]
  PIN rd_out[2051]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.665 0.070 791.735 ;
    END
  END rd_out[2051]
  PIN rd_out[2052]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.805 0.070 791.875 ;
    END
  END rd_out[2052]
  PIN rd_out[2053]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 791.945 0.070 792.015 ;
    END
  END rd_out[2053]
  PIN rd_out[2054]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.085 0.070 792.155 ;
    END
  END rd_out[2054]
  PIN rd_out[2055]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.225 0.070 792.295 ;
    END
  END rd_out[2055]
  PIN rd_out[2056]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.365 0.070 792.435 ;
    END
  END rd_out[2056]
  PIN rd_out[2057]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.505 0.070 792.575 ;
    END
  END rd_out[2057]
  PIN rd_out[2058]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.645 0.070 792.715 ;
    END
  END rd_out[2058]
  PIN rd_out[2059]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.785 0.070 792.855 ;
    END
  END rd_out[2059]
  PIN rd_out[2060]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 792.925 0.070 792.995 ;
    END
  END rd_out[2060]
  PIN rd_out[2061]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.065 0.070 793.135 ;
    END
  END rd_out[2061]
  PIN rd_out[2062]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.205 0.070 793.275 ;
    END
  END rd_out[2062]
  PIN rd_out[2063]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.345 0.070 793.415 ;
    END
  END rd_out[2063]
  PIN rd_out[2064]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.485 0.070 793.555 ;
    END
  END rd_out[2064]
  PIN rd_out[2065]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.625 0.070 793.695 ;
    END
  END rd_out[2065]
  PIN rd_out[2066]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.765 0.070 793.835 ;
    END
  END rd_out[2066]
  PIN rd_out[2067]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 793.905 0.070 793.975 ;
    END
  END rd_out[2067]
  PIN rd_out[2068]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.045 0.070 794.115 ;
    END
  END rd_out[2068]
  PIN rd_out[2069]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.185 0.070 794.255 ;
    END
  END rd_out[2069]
  PIN rd_out[2070]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.325 0.070 794.395 ;
    END
  END rd_out[2070]
  PIN rd_out[2071]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.465 0.070 794.535 ;
    END
  END rd_out[2071]
  PIN rd_out[2072]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.605 0.070 794.675 ;
    END
  END rd_out[2072]
  PIN rd_out[2073]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.745 0.070 794.815 ;
    END
  END rd_out[2073]
  PIN rd_out[2074]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 794.885 0.070 794.955 ;
    END
  END rd_out[2074]
  PIN rd_out[2075]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.025 0.070 795.095 ;
    END
  END rd_out[2075]
  PIN rd_out[2076]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.165 0.070 795.235 ;
    END
  END rd_out[2076]
  PIN rd_out[2077]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.305 0.070 795.375 ;
    END
  END rd_out[2077]
  PIN rd_out[2078]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.445 0.070 795.515 ;
    END
  END rd_out[2078]
  PIN rd_out[2079]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.585 0.070 795.655 ;
    END
  END rd_out[2079]
  PIN rd_out[2080]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.725 0.070 795.795 ;
    END
  END rd_out[2080]
  PIN rd_out[2081]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 795.865 0.070 795.935 ;
    END
  END rd_out[2081]
  PIN rd_out[2082]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.005 0.070 796.075 ;
    END
  END rd_out[2082]
  PIN rd_out[2083]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.145 0.070 796.215 ;
    END
  END rd_out[2083]
  PIN rd_out[2084]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.285 0.070 796.355 ;
    END
  END rd_out[2084]
  PIN rd_out[2085]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.425 0.070 796.495 ;
    END
  END rd_out[2085]
  PIN rd_out[2086]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.565 0.070 796.635 ;
    END
  END rd_out[2086]
  PIN rd_out[2087]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.705 0.070 796.775 ;
    END
  END rd_out[2087]
  PIN rd_out[2088]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.845 0.070 796.915 ;
    END
  END rd_out[2088]
  PIN rd_out[2089]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 796.985 0.070 797.055 ;
    END
  END rd_out[2089]
  PIN rd_out[2090]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.125 0.070 797.195 ;
    END
  END rd_out[2090]
  PIN rd_out[2091]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.265 0.070 797.335 ;
    END
  END rd_out[2091]
  PIN rd_out[2092]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.405 0.070 797.475 ;
    END
  END rd_out[2092]
  PIN rd_out[2093]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.545 0.070 797.615 ;
    END
  END rd_out[2093]
  PIN rd_out[2094]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.685 0.070 797.755 ;
    END
  END rd_out[2094]
  PIN rd_out[2095]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.825 0.070 797.895 ;
    END
  END rd_out[2095]
  PIN rd_out[2096]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 797.965 0.070 798.035 ;
    END
  END rd_out[2096]
  PIN rd_out[2097]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.105 0.070 798.175 ;
    END
  END rd_out[2097]
  PIN rd_out[2098]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.245 0.070 798.315 ;
    END
  END rd_out[2098]
  PIN rd_out[2099]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.385 0.070 798.455 ;
    END
  END rd_out[2099]
  PIN rd_out[2100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.525 0.070 798.595 ;
    END
  END rd_out[2100]
  PIN rd_out[2101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.665 0.070 798.735 ;
    END
  END rd_out[2101]
  PIN rd_out[2102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.805 0.070 798.875 ;
    END
  END rd_out[2102]
  PIN rd_out[2103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 798.945 0.070 799.015 ;
    END
  END rd_out[2103]
  PIN rd_out[2104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.085 0.070 799.155 ;
    END
  END rd_out[2104]
  PIN rd_out[2105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.225 0.070 799.295 ;
    END
  END rd_out[2105]
  PIN rd_out[2106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.365 0.070 799.435 ;
    END
  END rd_out[2106]
  PIN rd_out[2107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.505 0.070 799.575 ;
    END
  END rd_out[2107]
  PIN rd_out[2108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.645 0.070 799.715 ;
    END
  END rd_out[2108]
  PIN rd_out[2109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.785 0.070 799.855 ;
    END
  END rd_out[2109]
  PIN rd_out[2110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 799.925 0.070 799.995 ;
    END
  END rd_out[2110]
  PIN rd_out[2111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.065 0.070 800.135 ;
    END
  END rd_out[2111]
  PIN rd_out[2112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.205 0.070 800.275 ;
    END
  END rd_out[2112]
  PIN rd_out[2113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.345 0.070 800.415 ;
    END
  END rd_out[2113]
  PIN rd_out[2114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.485 0.070 800.555 ;
    END
  END rd_out[2114]
  PIN rd_out[2115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.625 0.070 800.695 ;
    END
  END rd_out[2115]
  PIN rd_out[2116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.765 0.070 800.835 ;
    END
  END rd_out[2116]
  PIN rd_out[2117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 800.905 0.070 800.975 ;
    END
  END rd_out[2117]
  PIN rd_out[2118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.045 0.070 801.115 ;
    END
  END rd_out[2118]
  PIN rd_out[2119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.185 0.070 801.255 ;
    END
  END rd_out[2119]
  PIN rd_out[2120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.325 0.070 801.395 ;
    END
  END rd_out[2120]
  PIN rd_out[2121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.465 0.070 801.535 ;
    END
  END rd_out[2121]
  PIN rd_out[2122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.605 0.070 801.675 ;
    END
  END rd_out[2122]
  PIN rd_out[2123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.745 0.070 801.815 ;
    END
  END rd_out[2123]
  PIN rd_out[2124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 801.885 0.070 801.955 ;
    END
  END rd_out[2124]
  PIN rd_out[2125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 802.025 0.070 802.095 ;
    END
  END rd_out[2125]
  PIN rd_out[2126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 802.165 0.070 802.235 ;
    END
  END rd_out[2126]
  PIN rd_out[2127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 802.305 0.070 802.375 ;
    END
  END rd_out[2127]
  PIN rd_out[2128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 802.445 0.070 802.515 ;
    END
  END rd_out[2128]
  PIN rd_out[2129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 802.585 0.070 802.655 ;
    END
  END rd_out[2129]
  PIN rd_out[2130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 802.725 0.070 802.795 ;
    END
  END rd_out[2130]
  PIN rd_out[2131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 802.865 0.070 802.935 ;
    END
  END rd_out[2131]
  PIN rd_out[2132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.005 0.070 803.075 ;
    END
  END rd_out[2132]
  PIN rd_out[2133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.145 0.070 803.215 ;
    END
  END rd_out[2133]
  PIN rd_out[2134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.285 0.070 803.355 ;
    END
  END rd_out[2134]
  PIN rd_out[2135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.425 0.070 803.495 ;
    END
  END rd_out[2135]
  PIN rd_out[2136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.565 0.070 803.635 ;
    END
  END rd_out[2136]
  PIN rd_out[2137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.705 0.070 803.775 ;
    END
  END rd_out[2137]
  PIN rd_out[2138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.845 0.070 803.915 ;
    END
  END rd_out[2138]
  PIN rd_out[2139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 803.985 0.070 804.055 ;
    END
  END rd_out[2139]
  PIN rd_out[2140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.125 0.070 804.195 ;
    END
  END rd_out[2140]
  PIN rd_out[2141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.265 0.070 804.335 ;
    END
  END rd_out[2141]
  PIN rd_out[2142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.405 0.070 804.475 ;
    END
  END rd_out[2142]
  PIN rd_out[2143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.545 0.070 804.615 ;
    END
  END rd_out[2143]
  PIN rd_out[2144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.685 0.070 804.755 ;
    END
  END rd_out[2144]
  PIN rd_out[2145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.825 0.070 804.895 ;
    END
  END rd_out[2145]
  PIN rd_out[2146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 804.965 0.070 805.035 ;
    END
  END rd_out[2146]
  PIN rd_out[2147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.105 0.070 805.175 ;
    END
  END rd_out[2147]
  PIN rd_out[2148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.245 0.070 805.315 ;
    END
  END rd_out[2148]
  PIN rd_out[2149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.385 0.070 805.455 ;
    END
  END rd_out[2149]
  PIN rd_out[2150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.525 0.070 805.595 ;
    END
  END rd_out[2150]
  PIN rd_out[2151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.665 0.070 805.735 ;
    END
  END rd_out[2151]
  PIN rd_out[2152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.805 0.070 805.875 ;
    END
  END rd_out[2152]
  PIN rd_out[2153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 805.945 0.070 806.015 ;
    END
  END rd_out[2153]
  PIN rd_out[2154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.085 0.070 806.155 ;
    END
  END rd_out[2154]
  PIN rd_out[2155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.225 0.070 806.295 ;
    END
  END rd_out[2155]
  PIN rd_out[2156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.365 0.070 806.435 ;
    END
  END rd_out[2156]
  PIN rd_out[2157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.505 0.070 806.575 ;
    END
  END rd_out[2157]
  PIN rd_out[2158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.645 0.070 806.715 ;
    END
  END rd_out[2158]
  PIN rd_out[2159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.785 0.070 806.855 ;
    END
  END rd_out[2159]
  PIN rd_out[2160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 806.925 0.070 806.995 ;
    END
  END rd_out[2160]
  PIN rd_out[2161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 807.065 0.070 807.135 ;
    END
  END rd_out[2161]
  PIN rd_out[2162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 807.205 0.070 807.275 ;
    END
  END rd_out[2162]
  PIN rd_out[2163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 807.345 0.070 807.415 ;
    END
  END rd_out[2163]
  PIN rd_out[2164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 807.485 0.070 807.555 ;
    END
  END rd_out[2164]
  PIN rd_out[2165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 807.625 0.070 807.695 ;
    END
  END rd_out[2165]
  PIN rd_out[2166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 807.765 0.070 807.835 ;
    END
  END rd_out[2166]
  PIN rd_out[2167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 807.905 0.070 807.975 ;
    END
  END rd_out[2167]
  PIN rd_out[2168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.045 0.070 808.115 ;
    END
  END rd_out[2168]
  PIN rd_out[2169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.185 0.070 808.255 ;
    END
  END rd_out[2169]
  PIN rd_out[2170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.325 0.070 808.395 ;
    END
  END rd_out[2170]
  PIN rd_out[2171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.465 0.070 808.535 ;
    END
  END rd_out[2171]
  PIN rd_out[2172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.605 0.070 808.675 ;
    END
  END rd_out[2172]
  PIN rd_out[2173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.745 0.070 808.815 ;
    END
  END rd_out[2173]
  PIN rd_out[2174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 808.885 0.070 808.955 ;
    END
  END rd_out[2174]
  PIN rd_out[2175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.025 0.070 809.095 ;
    END
  END rd_out[2175]
  PIN rd_out[2176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.165 0.070 809.235 ;
    END
  END rd_out[2176]
  PIN rd_out[2177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.305 0.070 809.375 ;
    END
  END rd_out[2177]
  PIN rd_out[2178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.445 0.070 809.515 ;
    END
  END rd_out[2178]
  PIN rd_out[2179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.585 0.070 809.655 ;
    END
  END rd_out[2179]
  PIN rd_out[2180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.725 0.070 809.795 ;
    END
  END rd_out[2180]
  PIN rd_out[2181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 809.865 0.070 809.935 ;
    END
  END rd_out[2181]
  PIN rd_out[2182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.005 0.070 810.075 ;
    END
  END rd_out[2182]
  PIN rd_out[2183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.145 0.070 810.215 ;
    END
  END rd_out[2183]
  PIN rd_out[2184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.285 0.070 810.355 ;
    END
  END rd_out[2184]
  PIN rd_out[2185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.425 0.070 810.495 ;
    END
  END rd_out[2185]
  PIN rd_out[2186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.565 0.070 810.635 ;
    END
  END rd_out[2186]
  PIN rd_out[2187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.705 0.070 810.775 ;
    END
  END rd_out[2187]
  PIN rd_out[2188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.845 0.070 810.915 ;
    END
  END rd_out[2188]
  PIN rd_out[2189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 810.985 0.070 811.055 ;
    END
  END rd_out[2189]
  PIN rd_out[2190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.125 0.070 811.195 ;
    END
  END rd_out[2190]
  PIN rd_out[2191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.265 0.070 811.335 ;
    END
  END rd_out[2191]
  PIN rd_out[2192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.405 0.070 811.475 ;
    END
  END rd_out[2192]
  PIN rd_out[2193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.545 0.070 811.615 ;
    END
  END rd_out[2193]
  PIN rd_out[2194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.685 0.070 811.755 ;
    END
  END rd_out[2194]
  PIN rd_out[2195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.825 0.070 811.895 ;
    END
  END rd_out[2195]
  PIN rd_out[2196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 811.965 0.070 812.035 ;
    END
  END rd_out[2196]
  PIN rd_out[2197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.105 0.070 812.175 ;
    END
  END rd_out[2197]
  PIN rd_out[2198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.245 0.070 812.315 ;
    END
  END rd_out[2198]
  PIN rd_out[2199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.385 0.070 812.455 ;
    END
  END rd_out[2199]
  PIN rd_out[2200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.525 0.070 812.595 ;
    END
  END rd_out[2200]
  PIN rd_out[2201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.665 0.070 812.735 ;
    END
  END rd_out[2201]
  PIN rd_out[2202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.805 0.070 812.875 ;
    END
  END rd_out[2202]
  PIN rd_out[2203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 812.945 0.070 813.015 ;
    END
  END rd_out[2203]
  PIN rd_out[2204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.085 0.070 813.155 ;
    END
  END rd_out[2204]
  PIN rd_out[2205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.225 0.070 813.295 ;
    END
  END rd_out[2205]
  PIN rd_out[2206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.365 0.070 813.435 ;
    END
  END rd_out[2206]
  PIN rd_out[2207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.505 0.070 813.575 ;
    END
  END rd_out[2207]
  PIN rd_out[2208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.645 0.070 813.715 ;
    END
  END rd_out[2208]
  PIN rd_out[2209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.785 0.070 813.855 ;
    END
  END rd_out[2209]
  PIN rd_out[2210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 813.925 0.070 813.995 ;
    END
  END rd_out[2210]
  PIN rd_out[2211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.065 0.070 814.135 ;
    END
  END rd_out[2211]
  PIN rd_out[2212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.205 0.070 814.275 ;
    END
  END rd_out[2212]
  PIN rd_out[2213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.345 0.070 814.415 ;
    END
  END rd_out[2213]
  PIN rd_out[2214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.485 0.070 814.555 ;
    END
  END rd_out[2214]
  PIN rd_out[2215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.625 0.070 814.695 ;
    END
  END rd_out[2215]
  PIN rd_out[2216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.765 0.070 814.835 ;
    END
  END rd_out[2216]
  PIN rd_out[2217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 814.905 0.070 814.975 ;
    END
  END rd_out[2217]
  PIN rd_out[2218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.045 0.070 815.115 ;
    END
  END rd_out[2218]
  PIN rd_out[2219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.185 0.070 815.255 ;
    END
  END rd_out[2219]
  PIN rd_out[2220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.325 0.070 815.395 ;
    END
  END rd_out[2220]
  PIN rd_out[2221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.465 0.070 815.535 ;
    END
  END rd_out[2221]
  PIN rd_out[2222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.605 0.070 815.675 ;
    END
  END rd_out[2222]
  PIN rd_out[2223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.745 0.070 815.815 ;
    END
  END rd_out[2223]
  PIN rd_out[2224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 815.885 0.070 815.955 ;
    END
  END rd_out[2224]
  PIN rd_out[2225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.025 0.070 816.095 ;
    END
  END rd_out[2225]
  PIN rd_out[2226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.165 0.070 816.235 ;
    END
  END rd_out[2226]
  PIN rd_out[2227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.305 0.070 816.375 ;
    END
  END rd_out[2227]
  PIN rd_out[2228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.445 0.070 816.515 ;
    END
  END rd_out[2228]
  PIN rd_out[2229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.585 0.070 816.655 ;
    END
  END rd_out[2229]
  PIN rd_out[2230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.725 0.070 816.795 ;
    END
  END rd_out[2230]
  PIN rd_out[2231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 816.865 0.070 816.935 ;
    END
  END rd_out[2231]
  PIN rd_out[2232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.005 0.070 817.075 ;
    END
  END rd_out[2232]
  PIN rd_out[2233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.145 0.070 817.215 ;
    END
  END rd_out[2233]
  PIN rd_out[2234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.285 0.070 817.355 ;
    END
  END rd_out[2234]
  PIN rd_out[2235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.425 0.070 817.495 ;
    END
  END rd_out[2235]
  PIN rd_out[2236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.565 0.070 817.635 ;
    END
  END rd_out[2236]
  PIN rd_out[2237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.705 0.070 817.775 ;
    END
  END rd_out[2237]
  PIN rd_out[2238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.845 0.070 817.915 ;
    END
  END rd_out[2238]
  PIN rd_out[2239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 817.985 0.070 818.055 ;
    END
  END rd_out[2239]
  PIN rd_out[2240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.125 0.070 818.195 ;
    END
  END rd_out[2240]
  PIN rd_out[2241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.265 0.070 818.335 ;
    END
  END rd_out[2241]
  PIN rd_out[2242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.405 0.070 818.475 ;
    END
  END rd_out[2242]
  PIN rd_out[2243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.545 0.070 818.615 ;
    END
  END rd_out[2243]
  PIN rd_out[2244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.685 0.070 818.755 ;
    END
  END rd_out[2244]
  PIN rd_out[2245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.825 0.070 818.895 ;
    END
  END rd_out[2245]
  PIN rd_out[2246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 818.965 0.070 819.035 ;
    END
  END rd_out[2246]
  PIN rd_out[2247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.105 0.070 819.175 ;
    END
  END rd_out[2247]
  PIN rd_out[2248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.245 0.070 819.315 ;
    END
  END rd_out[2248]
  PIN rd_out[2249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.385 0.070 819.455 ;
    END
  END rd_out[2249]
  PIN rd_out[2250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.525 0.070 819.595 ;
    END
  END rd_out[2250]
  PIN rd_out[2251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.665 0.070 819.735 ;
    END
  END rd_out[2251]
  PIN rd_out[2252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.805 0.070 819.875 ;
    END
  END rd_out[2252]
  PIN rd_out[2253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 819.945 0.070 820.015 ;
    END
  END rd_out[2253]
  PIN rd_out[2254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.085 0.070 820.155 ;
    END
  END rd_out[2254]
  PIN rd_out[2255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.225 0.070 820.295 ;
    END
  END rd_out[2255]
  PIN rd_out[2256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.365 0.070 820.435 ;
    END
  END rd_out[2256]
  PIN rd_out[2257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.505 0.070 820.575 ;
    END
  END rd_out[2257]
  PIN rd_out[2258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.645 0.070 820.715 ;
    END
  END rd_out[2258]
  PIN rd_out[2259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.785 0.070 820.855 ;
    END
  END rd_out[2259]
  PIN rd_out[2260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 820.925 0.070 820.995 ;
    END
  END rd_out[2260]
  PIN rd_out[2261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.065 0.070 821.135 ;
    END
  END rd_out[2261]
  PIN rd_out[2262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.205 0.070 821.275 ;
    END
  END rd_out[2262]
  PIN rd_out[2263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.345 0.070 821.415 ;
    END
  END rd_out[2263]
  PIN rd_out[2264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.485 0.070 821.555 ;
    END
  END rd_out[2264]
  PIN rd_out[2265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.625 0.070 821.695 ;
    END
  END rd_out[2265]
  PIN rd_out[2266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.765 0.070 821.835 ;
    END
  END rd_out[2266]
  PIN rd_out[2267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 821.905 0.070 821.975 ;
    END
  END rd_out[2267]
  PIN rd_out[2268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.045 0.070 822.115 ;
    END
  END rd_out[2268]
  PIN rd_out[2269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.185 0.070 822.255 ;
    END
  END rd_out[2269]
  PIN rd_out[2270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.325 0.070 822.395 ;
    END
  END rd_out[2270]
  PIN rd_out[2271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.465 0.070 822.535 ;
    END
  END rd_out[2271]
  PIN rd_out[2272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.605 0.070 822.675 ;
    END
  END rd_out[2272]
  PIN rd_out[2273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.745 0.070 822.815 ;
    END
  END rd_out[2273]
  PIN rd_out[2274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 822.885 0.070 822.955 ;
    END
  END rd_out[2274]
  PIN rd_out[2275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.025 0.070 823.095 ;
    END
  END rd_out[2275]
  PIN rd_out[2276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.165 0.070 823.235 ;
    END
  END rd_out[2276]
  PIN rd_out[2277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.305 0.070 823.375 ;
    END
  END rd_out[2277]
  PIN rd_out[2278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.445 0.070 823.515 ;
    END
  END rd_out[2278]
  PIN rd_out[2279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.585 0.070 823.655 ;
    END
  END rd_out[2279]
  PIN rd_out[2280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.725 0.070 823.795 ;
    END
  END rd_out[2280]
  PIN rd_out[2281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 823.865 0.070 823.935 ;
    END
  END rd_out[2281]
  PIN rd_out[2282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.005 0.070 824.075 ;
    END
  END rd_out[2282]
  PIN rd_out[2283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.145 0.070 824.215 ;
    END
  END rd_out[2283]
  PIN rd_out[2284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.285 0.070 824.355 ;
    END
  END rd_out[2284]
  PIN rd_out[2285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.425 0.070 824.495 ;
    END
  END rd_out[2285]
  PIN rd_out[2286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.565 0.070 824.635 ;
    END
  END rd_out[2286]
  PIN rd_out[2287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.705 0.070 824.775 ;
    END
  END rd_out[2287]
  PIN rd_out[2288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.845 0.070 824.915 ;
    END
  END rd_out[2288]
  PIN rd_out[2289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 824.985 0.070 825.055 ;
    END
  END rd_out[2289]
  PIN rd_out[2290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.125 0.070 825.195 ;
    END
  END rd_out[2290]
  PIN rd_out[2291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.265 0.070 825.335 ;
    END
  END rd_out[2291]
  PIN rd_out[2292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.405 0.070 825.475 ;
    END
  END rd_out[2292]
  PIN rd_out[2293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.545 0.070 825.615 ;
    END
  END rd_out[2293]
  PIN rd_out[2294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.685 0.070 825.755 ;
    END
  END rd_out[2294]
  PIN rd_out[2295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.825 0.070 825.895 ;
    END
  END rd_out[2295]
  PIN rd_out[2296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 825.965 0.070 826.035 ;
    END
  END rd_out[2296]
  PIN rd_out[2297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.105 0.070 826.175 ;
    END
  END rd_out[2297]
  PIN rd_out[2298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.245 0.070 826.315 ;
    END
  END rd_out[2298]
  PIN rd_out[2299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.385 0.070 826.455 ;
    END
  END rd_out[2299]
  PIN rd_out[2300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.525 0.070 826.595 ;
    END
  END rd_out[2300]
  PIN rd_out[2301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.665 0.070 826.735 ;
    END
  END rd_out[2301]
  PIN rd_out[2302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.805 0.070 826.875 ;
    END
  END rd_out[2302]
  PIN rd_out[2303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 826.945 0.070 827.015 ;
    END
  END rd_out[2303]
  PIN rd_out[2304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.085 0.070 827.155 ;
    END
  END rd_out[2304]
  PIN rd_out[2305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.225 0.070 827.295 ;
    END
  END rd_out[2305]
  PIN rd_out[2306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.365 0.070 827.435 ;
    END
  END rd_out[2306]
  PIN rd_out[2307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.505 0.070 827.575 ;
    END
  END rd_out[2307]
  PIN rd_out[2308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.645 0.070 827.715 ;
    END
  END rd_out[2308]
  PIN rd_out[2309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.785 0.070 827.855 ;
    END
  END rd_out[2309]
  PIN rd_out[2310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 827.925 0.070 827.995 ;
    END
  END rd_out[2310]
  PIN rd_out[2311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.065 0.070 828.135 ;
    END
  END rd_out[2311]
  PIN rd_out[2312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.205 0.070 828.275 ;
    END
  END rd_out[2312]
  PIN rd_out[2313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.345 0.070 828.415 ;
    END
  END rd_out[2313]
  PIN rd_out[2314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.485 0.070 828.555 ;
    END
  END rd_out[2314]
  PIN rd_out[2315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.625 0.070 828.695 ;
    END
  END rd_out[2315]
  PIN rd_out[2316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.765 0.070 828.835 ;
    END
  END rd_out[2316]
  PIN rd_out[2317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 828.905 0.070 828.975 ;
    END
  END rd_out[2317]
  PIN rd_out[2318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.045 0.070 829.115 ;
    END
  END rd_out[2318]
  PIN rd_out[2319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.185 0.070 829.255 ;
    END
  END rd_out[2319]
  PIN rd_out[2320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.325 0.070 829.395 ;
    END
  END rd_out[2320]
  PIN rd_out[2321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.465 0.070 829.535 ;
    END
  END rd_out[2321]
  PIN rd_out[2322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.605 0.070 829.675 ;
    END
  END rd_out[2322]
  PIN rd_out[2323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.745 0.070 829.815 ;
    END
  END rd_out[2323]
  PIN rd_out[2324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 829.885 0.070 829.955 ;
    END
  END rd_out[2324]
  PIN rd_out[2325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.025 0.070 830.095 ;
    END
  END rd_out[2325]
  PIN rd_out[2326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.165 0.070 830.235 ;
    END
  END rd_out[2326]
  PIN rd_out[2327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.305 0.070 830.375 ;
    END
  END rd_out[2327]
  PIN rd_out[2328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.445 0.070 830.515 ;
    END
  END rd_out[2328]
  PIN rd_out[2329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.585 0.070 830.655 ;
    END
  END rd_out[2329]
  PIN rd_out[2330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.725 0.070 830.795 ;
    END
  END rd_out[2330]
  PIN rd_out[2331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 830.865 0.070 830.935 ;
    END
  END rd_out[2331]
  PIN rd_out[2332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.005 0.070 831.075 ;
    END
  END rd_out[2332]
  PIN rd_out[2333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.145 0.070 831.215 ;
    END
  END rd_out[2333]
  PIN rd_out[2334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.285 0.070 831.355 ;
    END
  END rd_out[2334]
  PIN rd_out[2335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.425 0.070 831.495 ;
    END
  END rd_out[2335]
  PIN rd_out[2336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.565 0.070 831.635 ;
    END
  END rd_out[2336]
  PIN rd_out[2337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.705 0.070 831.775 ;
    END
  END rd_out[2337]
  PIN rd_out[2338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.845 0.070 831.915 ;
    END
  END rd_out[2338]
  PIN rd_out[2339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 831.985 0.070 832.055 ;
    END
  END rd_out[2339]
  PIN rd_out[2340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.125 0.070 832.195 ;
    END
  END rd_out[2340]
  PIN rd_out[2341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.265 0.070 832.335 ;
    END
  END rd_out[2341]
  PIN rd_out[2342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.405 0.070 832.475 ;
    END
  END rd_out[2342]
  PIN rd_out[2343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.545 0.070 832.615 ;
    END
  END rd_out[2343]
  PIN rd_out[2344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.685 0.070 832.755 ;
    END
  END rd_out[2344]
  PIN rd_out[2345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.825 0.070 832.895 ;
    END
  END rd_out[2345]
  PIN rd_out[2346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 832.965 0.070 833.035 ;
    END
  END rd_out[2346]
  PIN rd_out[2347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.105 0.070 833.175 ;
    END
  END rd_out[2347]
  PIN rd_out[2348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.245 0.070 833.315 ;
    END
  END rd_out[2348]
  PIN rd_out[2349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.385 0.070 833.455 ;
    END
  END rd_out[2349]
  PIN rd_out[2350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.525 0.070 833.595 ;
    END
  END rd_out[2350]
  PIN rd_out[2351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.665 0.070 833.735 ;
    END
  END rd_out[2351]
  PIN rd_out[2352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.805 0.070 833.875 ;
    END
  END rd_out[2352]
  PIN rd_out[2353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 833.945 0.070 834.015 ;
    END
  END rd_out[2353]
  PIN rd_out[2354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.085 0.070 834.155 ;
    END
  END rd_out[2354]
  PIN rd_out[2355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.225 0.070 834.295 ;
    END
  END rd_out[2355]
  PIN rd_out[2356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.365 0.070 834.435 ;
    END
  END rd_out[2356]
  PIN rd_out[2357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.505 0.070 834.575 ;
    END
  END rd_out[2357]
  PIN rd_out[2358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.645 0.070 834.715 ;
    END
  END rd_out[2358]
  PIN rd_out[2359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.785 0.070 834.855 ;
    END
  END rd_out[2359]
  PIN rd_out[2360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 834.925 0.070 834.995 ;
    END
  END rd_out[2360]
  PIN rd_out[2361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.065 0.070 835.135 ;
    END
  END rd_out[2361]
  PIN rd_out[2362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.205 0.070 835.275 ;
    END
  END rd_out[2362]
  PIN rd_out[2363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.345 0.070 835.415 ;
    END
  END rd_out[2363]
  PIN rd_out[2364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.485 0.070 835.555 ;
    END
  END rd_out[2364]
  PIN rd_out[2365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.625 0.070 835.695 ;
    END
  END rd_out[2365]
  PIN rd_out[2366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.765 0.070 835.835 ;
    END
  END rd_out[2366]
  PIN rd_out[2367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 835.905 0.070 835.975 ;
    END
  END rd_out[2367]
  PIN rd_out[2368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.045 0.070 836.115 ;
    END
  END rd_out[2368]
  PIN rd_out[2369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.185 0.070 836.255 ;
    END
  END rd_out[2369]
  PIN rd_out[2370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.325 0.070 836.395 ;
    END
  END rd_out[2370]
  PIN rd_out[2371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.465 0.070 836.535 ;
    END
  END rd_out[2371]
  PIN rd_out[2372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.605 0.070 836.675 ;
    END
  END rd_out[2372]
  PIN rd_out[2373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.745 0.070 836.815 ;
    END
  END rd_out[2373]
  PIN rd_out[2374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 836.885 0.070 836.955 ;
    END
  END rd_out[2374]
  PIN rd_out[2375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.025 0.070 837.095 ;
    END
  END rd_out[2375]
  PIN rd_out[2376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.165 0.070 837.235 ;
    END
  END rd_out[2376]
  PIN rd_out[2377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.305 0.070 837.375 ;
    END
  END rd_out[2377]
  PIN rd_out[2378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.445 0.070 837.515 ;
    END
  END rd_out[2378]
  PIN rd_out[2379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.585 0.070 837.655 ;
    END
  END rd_out[2379]
  PIN rd_out[2380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.725 0.070 837.795 ;
    END
  END rd_out[2380]
  PIN rd_out[2381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 837.865 0.070 837.935 ;
    END
  END rd_out[2381]
  PIN rd_out[2382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.005 0.070 838.075 ;
    END
  END rd_out[2382]
  PIN rd_out[2383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.145 0.070 838.215 ;
    END
  END rd_out[2383]
  PIN rd_out[2384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.285 0.070 838.355 ;
    END
  END rd_out[2384]
  PIN rd_out[2385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.425 0.070 838.495 ;
    END
  END rd_out[2385]
  PIN rd_out[2386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.565 0.070 838.635 ;
    END
  END rd_out[2386]
  PIN rd_out[2387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.705 0.070 838.775 ;
    END
  END rd_out[2387]
  PIN rd_out[2388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.845 0.070 838.915 ;
    END
  END rd_out[2388]
  PIN rd_out[2389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 838.985 0.070 839.055 ;
    END
  END rd_out[2389]
  PIN rd_out[2390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.125 0.070 839.195 ;
    END
  END rd_out[2390]
  PIN rd_out[2391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.265 0.070 839.335 ;
    END
  END rd_out[2391]
  PIN rd_out[2392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.405 0.070 839.475 ;
    END
  END rd_out[2392]
  PIN rd_out[2393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.545 0.070 839.615 ;
    END
  END rd_out[2393]
  PIN rd_out[2394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.685 0.070 839.755 ;
    END
  END rd_out[2394]
  PIN rd_out[2395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.825 0.070 839.895 ;
    END
  END rd_out[2395]
  PIN rd_out[2396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 839.965 0.070 840.035 ;
    END
  END rd_out[2396]
  PIN rd_out[2397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.105 0.070 840.175 ;
    END
  END rd_out[2397]
  PIN rd_out[2398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.245 0.070 840.315 ;
    END
  END rd_out[2398]
  PIN rd_out[2399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.385 0.070 840.455 ;
    END
  END rd_out[2399]
  PIN rd_out[2400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.525 0.070 840.595 ;
    END
  END rd_out[2400]
  PIN rd_out[2401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.665 0.070 840.735 ;
    END
  END rd_out[2401]
  PIN rd_out[2402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.805 0.070 840.875 ;
    END
  END rd_out[2402]
  PIN rd_out[2403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 840.945 0.070 841.015 ;
    END
  END rd_out[2403]
  PIN rd_out[2404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.085 0.070 841.155 ;
    END
  END rd_out[2404]
  PIN rd_out[2405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.225 0.070 841.295 ;
    END
  END rd_out[2405]
  PIN rd_out[2406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.365 0.070 841.435 ;
    END
  END rd_out[2406]
  PIN rd_out[2407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.505 0.070 841.575 ;
    END
  END rd_out[2407]
  PIN rd_out[2408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.645 0.070 841.715 ;
    END
  END rd_out[2408]
  PIN rd_out[2409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.785 0.070 841.855 ;
    END
  END rd_out[2409]
  PIN rd_out[2410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 841.925 0.070 841.995 ;
    END
  END rd_out[2410]
  PIN rd_out[2411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.065 0.070 842.135 ;
    END
  END rd_out[2411]
  PIN rd_out[2412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.205 0.070 842.275 ;
    END
  END rd_out[2412]
  PIN rd_out[2413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.345 0.070 842.415 ;
    END
  END rd_out[2413]
  PIN rd_out[2414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.485 0.070 842.555 ;
    END
  END rd_out[2414]
  PIN rd_out[2415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.625 0.070 842.695 ;
    END
  END rd_out[2415]
  PIN rd_out[2416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.765 0.070 842.835 ;
    END
  END rd_out[2416]
  PIN rd_out[2417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 842.905 0.070 842.975 ;
    END
  END rd_out[2417]
  PIN rd_out[2418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.045 0.070 843.115 ;
    END
  END rd_out[2418]
  PIN rd_out[2419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.185 0.070 843.255 ;
    END
  END rd_out[2419]
  PIN rd_out[2420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.325 0.070 843.395 ;
    END
  END rd_out[2420]
  PIN rd_out[2421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.465 0.070 843.535 ;
    END
  END rd_out[2421]
  PIN rd_out[2422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.605 0.070 843.675 ;
    END
  END rd_out[2422]
  PIN rd_out[2423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.745 0.070 843.815 ;
    END
  END rd_out[2423]
  PIN rd_out[2424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 843.885 0.070 843.955 ;
    END
  END rd_out[2424]
  PIN rd_out[2425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.025 0.070 844.095 ;
    END
  END rd_out[2425]
  PIN rd_out[2426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.165 0.070 844.235 ;
    END
  END rd_out[2426]
  PIN rd_out[2427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.305 0.070 844.375 ;
    END
  END rd_out[2427]
  PIN rd_out[2428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.445 0.070 844.515 ;
    END
  END rd_out[2428]
  PIN rd_out[2429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.585 0.070 844.655 ;
    END
  END rd_out[2429]
  PIN rd_out[2430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.725 0.070 844.795 ;
    END
  END rd_out[2430]
  PIN rd_out[2431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 844.865 0.070 844.935 ;
    END
  END rd_out[2431]
  PIN rd_out[2432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.005 0.070 845.075 ;
    END
  END rd_out[2432]
  PIN rd_out[2433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.145 0.070 845.215 ;
    END
  END rd_out[2433]
  PIN rd_out[2434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.285 0.070 845.355 ;
    END
  END rd_out[2434]
  PIN rd_out[2435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.425 0.070 845.495 ;
    END
  END rd_out[2435]
  PIN rd_out[2436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.565 0.070 845.635 ;
    END
  END rd_out[2436]
  PIN rd_out[2437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.705 0.070 845.775 ;
    END
  END rd_out[2437]
  PIN rd_out[2438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.845 0.070 845.915 ;
    END
  END rd_out[2438]
  PIN rd_out[2439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 845.985 0.070 846.055 ;
    END
  END rd_out[2439]
  PIN rd_out[2440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.125 0.070 846.195 ;
    END
  END rd_out[2440]
  PIN rd_out[2441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.265 0.070 846.335 ;
    END
  END rd_out[2441]
  PIN rd_out[2442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.405 0.070 846.475 ;
    END
  END rd_out[2442]
  PIN rd_out[2443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.545 0.070 846.615 ;
    END
  END rd_out[2443]
  PIN rd_out[2444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.685 0.070 846.755 ;
    END
  END rd_out[2444]
  PIN rd_out[2445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.825 0.070 846.895 ;
    END
  END rd_out[2445]
  PIN rd_out[2446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 846.965 0.070 847.035 ;
    END
  END rd_out[2446]
  PIN rd_out[2447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.105 0.070 847.175 ;
    END
  END rd_out[2447]
  PIN rd_out[2448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.245 0.070 847.315 ;
    END
  END rd_out[2448]
  PIN rd_out[2449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.385 0.070 847.455 ;
    END
  END rd_out[2449]
  PIN rd_out[2450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.525 0.070 847.595 ;
    END
  END rd_out[2450]
  PIN rd_out[2451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.665 0.070 847.735 ;
    END
  END rd_out[2451]
  PIN rd_out[2452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.805 0.070 847.875 ;
    END
  END rd_out[2452]
  PIN rd_out[2453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 847.945 0.070 848.015 ;
    END
  END rd_out[2453]
  PIN rd_out[2454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.085 0.070 848.155 ;
    END
  END rd_out[2454]
  PIN rd_out[2455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.225 0.070 848.295 ;
    END
  END rd_out[2455]
  PIN rd_out[2456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.365 0.070 848.435 ;
    END
  END rd_out[2456]
  PIN rd_out[2457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.505 0.070 848.575 ;
    END
  END rd_out[2457]
  PIN rd_out[2458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.645 0.070 848.715 ;
    END
  END rd_out[2458]
  PIN rd_out[2459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.785 0.070 848.855 ;
    END
  END rd_out[2459]
  PIN rd_out[2460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 848.925 0.070 848.995 ;
    END
  END rd_out[2460]
  PIN rd_out[2461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.065 0.070 849.135 ;
    END
  END rd_out[2461]
  PIN rd_out[2462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.205 0.070 849.275 ;
    END
  END rd_out[2462]
  PIN rd_out[2463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.345 0.070 849.415 ;
    END
  END rd_out[2463]
  PIN rd_out[2464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.485 0.070 849.555 ;
    END
  END rd_out[2464]
  PIN rd_out[2465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.625 0.070 849.695 ;
    END
  END rd_out[2465]
  PIN rd_out[2466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.765 0.070 849.835 ;
    END
  END rd_out[2466]
  PIN rd_out[2467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 849.905 0.070 849.975 ;
    END
  END rd_out[2467]
  PIN rd_out[2468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.045 0.070 850.115 ;
    END
  END rd_out[2468]
  PIN rd_out[2469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.185 0.070 850.255 ;
    END
  END rd_out[2469]
  PIN rd_out[2470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.325 0.070 850.395 ;
    END
  END rd_out[2470]
  PIN rd_out[2471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.465 0.070 850.535 ;
    END
  END rd_out[2471]
  PIN rd_out[2472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.605 0.070 850.675 ;
    END
  END rd_out[2472]
  PIN rd_out[2473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.745 0.070 850.815 ;
    END
  END rd_out[2473]
  PIN rd_out[2474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 850.885 0.070 850.955 ;
    END
  END rd_out[2474]
  PIN rd_out[2475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.025 0.070 851.095 ;
    END
  END rd_out[2475]
  PIN rd_out[2476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.165 0.070 851.235 ;
    END
  END rd_out[2476]
  PIN rd_out[2477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.305 0.070 851.375 ;
    END
  END rd_out[2477]
  PIN rd_out[2478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.445 0.070 851.515 ;
    END
  END rd_out[2478]
  PIN rd_out[2479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.585 0.070 851.655 ;
    END
  END rd_out[2479]
  PIN rd_out[2480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.725 0.070 851.795 ;
    END
  END rd_out[2480]
  PIN rd_out[2481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 851.865 0.070 851.935 ;
    END
  END rd_out[2481]
  PIN rd_out[2482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.005 0.070 852.075 ;
    END
  END rd_out[2482]
  PIN rd_out[2483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.145 0.070 852.215 ;
    END
  END rd_out[2483]
  PIN rd_out[2484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.285 0.070 852.355 ;
    END
  END rd_out[2484]
  PIN rd_out[2485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.425 0.070 852.495 ;
    END
  END rd_out[2485]
  PIN rd_out[2486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.565 0.070 852.635 ;
    END
  END rd_out[2486]
  PIN rd_out[2487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.705 0.070 852.775 ;
    END
  END rd_out[2487]
  PIN rd_out[2488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.845 0.070 852.915 ;
    END
  END rd_out[2488]
  PIN rd_out[2489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 852.985 0.070 853.055 ;
    END
  END rd_out[2489]
  PIN rd_out[2490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.125 0.070 853.195 ;
    END
  END rd_out[2490]
  PIN rd_out[2491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.265 0.070 853.335 ;
    END
  END rd_out[2491]
  PIN rd_out[2492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.405 0.070 853.475 ;
    END
  END rd_out[2492]
  PIN rd_out[2493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.545 0.070 853.615 ;
    END
  END rd_out[2493]
  PIN rd_out[2494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.685 0.070 853.755 ;
    END
  END rd_out[2494]
  PIN rd_out[2495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.825 0.070 853.895 ;
    END
  END rd_out[2495]
  PIN rd_out[2496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 853.965 0.070 854.035 ;
    END
  END rd_out[2496]
  PIN rd_out[2497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.105 0.070 854.175 ;
    END
  END rd_out[2497]
  PIN rd_out[2498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.245 0.070 854.315 ;
    END
  END rd_out[2498]
  PIN rd_out[2499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.385 0.070 854.455 ;
    END
  END rd_out[2499]
  PIN rd_out[2500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.525 0.070 854.595 ;
    END
  END rd_out[2500]
  PIN rd_out[2501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.665 0.070 854.735 ;
    END
  END rd_out[2501]
  PIN rd_out[2502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.805 0.070 854.875 ;
    END
  END rd_out[2502]
  PIN rd_out[2503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 854.945 0.070 855.015 ;
    END
  END rd_out[2503]
  PIN rd_out[2504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.085 0.070 855.155 ;
    END
  END rd_out[2504]
  PIN rd_out[2505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.225 0.070 855.295 ;
    END
  END rd_out[2505]
  PIN rd_out[2506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.365 0.070 855.435 ;
    END
  END rd_out[2506]
  PIN rd_out[2507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.505 0.070 855.575 ;
    END
  END rd_out[2507]
  PIN rd_out[2508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.645 0.070 855.715 ;
    END
  END rd_out[2508]
  PIN rd_out[2509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.785 0.070 855.855 ;
    END
  END rd_out[2509]
  PIN rd_out[2510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 855.925 0.070 855.995 ;
    END
  END rd_out[2510]
  PIN rd_out[2511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.065 0.070 856.135 ;
    END
  END rd_out[2511]
  PIN rd_out[2512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.205 0.070 856.275 ;
    END
  END rd_out[2512]
  PIN rd_out[2513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.345 0.070 856.415 ;
    END
  END rd_out[2513]
  PIN rd_out[2514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.485 0.070 856.555 ;
    END
  END rd_out[2514]
  PIN rd_out[2515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.625 0.070 856.695 ;
    END
  END rd_out[2515]
  PIN rd_out[2516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.765 0.070 856.835 ;
    END
  END rd_out[2516]
  PIN rd_out[2517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 856.905 0.070 856.975 ;
    END
  END rd_out[2517]
  PIN rd_out[2518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.045 0.070 857.115 ;
    END
  END rd_out[2518]
  PIN rd_out[2519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.185 0.070 857.255 ;
    END
  END rd_out[2519]
  PIN rd_out[2520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.325 0.070 857.395 ;
    END
  END rd_out[2520]
  PIN rd_out[2521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.465 0.070 857.535 ;
    END
  END rd_out[2521]
  PIN rd_out[2522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.605 0.070 857.675 ;
    END
  END rd_out[2522]
  PIN rd_out[2523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.745 0.070 857.815 ;
    END
  END rd_out[2523]
  PIN rd_out[2524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 857.885 0.070 857.955 ;
    END
  END rd_out[2524]
  PIN rd_out[2525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.025 0.070 858.095 ;
    END
  END rd_out[2525]
  PIN rd_out[2526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.165 0.070 858.235 ;
    END
  END rd_out[2526]
  PIN rd_out[2527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.305 0.070 858.375 ;
    END
  END rd_out[2527]
  PIN rd_out[2528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.445 0.070 858.515 ;
    END
  END rd_out[2528]
  PIN rd_out[2529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.585 0.070 858.655 ;
    END
  END rd_out[2529]
  PIN rd_out[2530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.725 0.070 858.795 ;
    END
  END rd_out[2530]
  PIN rd_out[2531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 858.865 0.070 858.935 ;
    END
  END rd_out[2531]
  PIN rd_out[2532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.005 0.070 859.075 ;
    END
  END rd_out[2532]
  PIN rd_out[2533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.145 0.070 859.215 ;
    END
  END rd_out[2533]
  PIN rd_out[2534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.285 0.070 859.355 ;
    END
  END rd_out[2534]
  PIN rd_out[2535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.425 0.070 859.495 ;
    END
  END rd_out[2535]
  PIN rd_out[2536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.565 0.070 859.635 ;
    END
  END rd_out[2536]
  PIN rd_out[2537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.705 0.070 859.775 ;
    END
  END rd_out[2537]
  PIN rd_out[2538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.845 0.070 859.915 ;
    END
  END rd_out[2538]
  PIN rd_out[2539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 859.985 0.070 860.055 ;
    END
  END rd_out[2539]
  PIN rd_out[2540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.125 0.070 860.195 ;
    END
  END rd_out[2540]
  PIN rd_out[2541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.265 0.070 860.335 ;
    END
  END rd_out[2541]
  PIN rd_out[2542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.405 0.070 860.475 ;
    END
  END rd_out[2542]
  PIN rd_out[2543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.545 0.070 860.615 ;
    END
  END rd_out[2543]
  PIN rd_out[2544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.685 0.070 860.755 ;
    END
  END rd_out[2544]
  PIN rd_out[2545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.825 0.070 860.895 ;
    END
  END rd_out[2545]
  PIN rd_out[2546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 860.965 0.070 861.035 ;
    END
  END rd_out[2546]
  PIN rd_out[2547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.105 0.070 861.175 ;
    END
  END rd_out[2547]
  PIN rd_out[2548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.245 0.070 861.315 ;
    END
  END rd_out[2548]
  PIN rd_out[2549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.385 0.070 861.455 ;
    END
  END rd_out[2549]
  PIN rd_out[2550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.525 0.070 861.595 ;
    END
  END rd_out[2550]
  PIN rd_out[2551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.665 0.070 861.735 ;
    END
  END rd_out[2551]
  PIN rd_out[2552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.805 0.070 861.875 ;
    END
  END rd_out[2552]
  PIN rd_out[2553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 861.945 0.070 862.015 ;
    END
  END rd_out[2553]
  PIN rd_out[2554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.085 0.070 862.155 ;
    END
  END rd_out[2554]
  PIN rd_out[2555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.225 0.070 862.295 ;
    END
  END rd_out[2555]
  PIN rd_out[2556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.365 0.070 862.435 ;
    END
  END rd_out[2556]
  PIN rd_out[2557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.505 0.070 862.575 ;
    END
  END rd_out[2557]
  PIN rd_out[2558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.645 0.070 862.715 ;
    END
  END rd_out[2558]
  PIN rd_out[2559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.785 0.070 862.855 ;
    END
  END rd_out[2559]
  PIN rd_out[2560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 862.925 0.070 862.995 ;
    END
  END rd_out[2560]
  PIN rd_out[2561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.065 0.070 863.135 ;
    END
  END rd_out[2561]
  PIN rd_out[2562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.205 0.070 863.275 ;
    END
  END rd_out[2562]
  PIN rd_out[2563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.345 0.070 863.415 ;
    END
  END rd_out[2563]
  PIN rd_out[2564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.485 0.070 863.555 ;
    END
  END rd_out[2564]
  PIN rd_out[2565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.625 0.070 863.695 ;
    END
  END rd_out[2565]
  PIN rd_out[2566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.765 0.070 863.835 ;
    END
  END rd_out[2566]
  PIN rd_out[2567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 863.905 0.070 863.975 ;
    END
  END rd_out[2567]
  PIN rd_out[2568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.045 0.070 864.115 ;
    END
  END rd_out[2568]
  PIN rd_out[2569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.185 0.070 864.255 ;
    END
  END rd_out[2569]
  PIN rd_out[2570]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.325 0.070 864.395 ;
    END
  END rd_out[2570]
  PIN rd_out[2571]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.465 0.070 864.535 ;
    END
  END rd_out[2571]
  PIN rd_out[2572]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.605 0.070 864.675 ;
    END
  END rd_out[2572]
  PIN rd_out[2573]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.745 0.070 864.815 ;
    END
  END rd_out[2573]
  PIN rd_out[2574]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 864.885 0.070 864.955 ;
    END
  END rd_out[2574]
  PIN rd_out[2575]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.025 0.070 865.095 ;
    END
  END rd_out[2575]
  PIN rd_out[2576]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.165 0.070 865.235 ;
    END
  END rd_out[2576]
  PIN rd_out[2577]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.305 0.070 865.375 ;
    END
  END rd_out[2577]
  PIN rd_out[2578]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.445 0.070 865.515 ;
    END
  END rd_out[2578]
  PIN rd_out[2579]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.585 0.070 865.655 ;
    END
  END rd_out[2579]
  PIN rd_out[2580]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.725 0.070 865.795 ;
    END
  END rd_out[2580]
  PIN rd_out[2581]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 865.865 0.070 865.935 ;
    END
  END rd_out[2581]
  PIN rd_out[2582]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.005 0.070 866.075 ;
    END
  END rd_out[2582]
  PIN rd_out[2583]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.145 0.070 866.215 ;
    END
  END rd_out[2583]
  PIN rd_out[2584]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.285 0.070 866.355 ;
    END
  END rd_out[2584]
  PIN rd_out[2585]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.425 0.070 866.495 ;
    END
  END rd_out[2585]
  PIN rd_out[2586]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.565 0.070 866.635 ;
    END
  END rd_out[2586]
  PIN rd_out[2587]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.705 0.070 866.775 ;
    END
  END rd_out[2587]
  PIN rd_out[2588]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.845 0.070 866.915 ;
    END
  END rd_out[2588]
  PIN rd_out[2589]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 866.985 0.070 867.055 ;
    END
  END rd_out[2589]
  PIN rd_out[2590]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.125 0.070 867.195 ;
    END
  END rd_out[2590]
  PIN rd_out[2591]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.265 0.070 867.335 ;
    END
  END rd_out[2591]
  PIN rd_out[2592]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.405 0.070 867.475 ;
    END
  END rd_out[2592]
  PIN rd_out[2593]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.545 0.070 867.615 ;
    END
  END rd_out[2593]
  PIN rd_out[2594]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.685 0.070 867.755 ;
    END
  END rd_out[2594]
  PIN rd_out[2595]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.825 0.070 867.895 ;
    END
  END rd_out[2595]
  PIN rd_out[2596]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 867.965 0.070 868.035 ;
    END
  END rd_out[2596]
  PIN rd_out[2597]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.105 0.070 868.175 ;
    END
  END rd_out[2597]
  PIN rd_out[2598]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.245 0.070 868.315 ;
    END
  END rd_out[2598]
  PIN rd_out[2599]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.385 0.070 868.455 ;
    END
  END rd_out[2599]
  PIN rd_out[2600]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.525 0.070 868.595 ;
    END
  END rd_out[2600]
  PIN rd_out[2601]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.665 0.070 868.735 ;
    END
  END rd_out[2601]
  PIN rd_out[2602]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.805 0.070 868.875 ;
    END
  END rd_out[2602]
  PIN rd_out[2603]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 868.945 0.070 869.015 ;
    END
  END rd_out[2603]
  PIN rd_out[2604]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.085 0.070 869.155 ;
    END
  END rd_out[2604]
  PIN rd_out[2605]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.225 0.070 869.295 ;
    END
  END rd_out[2605]
  PIN rd_out[2606]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.365 0.070 869.435 ;
    END
  END rd_out[2606]
  PIN rd_out[2607]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.505 0.070 869.575 ;
    END
  END rd_out[2607]
  PIN rd_out[2608]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.645 0.070 869.715 ;
    END
  END rd_out[2608]
  PIN rd_out[2609]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.785 0.070 869.855 ;
    END
  END rd_out[2609]
  PIN rd_out[2610]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 869.925 0.070 869.995 ;
    END
  END rd_out[2610]
  PIN rd_out[2611]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.065 0.070 870.135 ;
    END
  END rd_out[2611]
  PIN rd_out[2612]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.205 0.070 870.275 ;
    END
  END rd_out[2612]
  PIN rd_out[2613]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.345 0.070 870.415 ;
    END
  END rd_out[2613]
  PIN rd_out[2614]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.485 0.070 870.555 ;
    END
  END rd_out[2614]
  PIN rd_out[2615]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.625 0.070 870.695 ;
    END
  END rd_out[2615]
  PIN rd_out[2616]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.765 0.070 870.835 ;
    END
  END rd_out[2616]
  PIN rd_out[2617]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 870.905 0.070 870.975 ;
    END
  END rd_out[2617]
  PIN rd_out[2618]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.045 0.070 871.115 ;
    END
  END rd_out[2618]
  PIN rd_out[2619]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.185 0.070 871.255 ;
    END
  END rd_out[2619]
  PIN rd_out[2620]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.325 0.070 871.395 ;
    END
  END rd_out[2620]
  PIN rd_out[2621]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.465 0.070 871.535 ;
    END
  END rd_out[2621]
  PIN rd_out[2622]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.605 0.070 871.675 ;
    END
  END rd_out[2622]
  PIN rd_out[2623]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.745 0.070 871.815 ;
    END
  END rd_out[2623]
  PIN rd_out[2624]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 871.885 0.070 871.955 ;
    END
  END rd_out[2624]
  PIN rd_out[2625]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.025 0.070 872.095 ;
    END
  END rd_out[2625]
  PIN rd_out[2626]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.165 0.070 872.235 ;
    END
  END rd_out[2626]
  PIN rd_out[2627]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.305 0.070 872.375 ;
    END
  END rd_out[2627]
  PIN rd_out[2628]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.445 0.070 872.515 ;
    END
  END rd_out[2628]
  PIN rd_out[2629]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.585 0.070 872.655 ;
    END
  END rd_out[2629]
  PIN rd_out[2630]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.725 0.070 872.795 ;
    END
  END rd_out[2630]
  PIN rd_out[2631]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 872.865 0.070 872.935 ;
    END
  END rd_out[2631]
  PIN rd_out[2632]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.005 0.070 873.075 ;
    END
  END rd_out[2632]
  PIN rd_out[2633]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.145 0.070 873.215 ;
    END
  END rd_out[2633]
  PIN rd_out[2634]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.285 0.070 873.355 ;
    END
  END rd_out[2634]
  PIN rd_out[2635]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.425 0.070 873.495 ;
    END
  END rd_out[2635]
  PIN rd_out[2636]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.565 0.070 873.635 ;
    END
  END rd_out[2636]
  PIN rd_out[2637]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.705 0.070 873.775 ;
    END
  END rd_out[2637]
  PIN rd_out[2638]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.845 0.070 873.915 ;
    END
  END rd_out[2638]
  PIN rd_out[2639]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 873.985 0.070 874.055 ;
    END
  END rd_out[2639]
  PIN rd_out[2640]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.125 0.070 874.195 ;
    END
  END rd_out[2640]
  PIN rd_out[2641]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.265 0.070 874.335 ;
    END
  END rd_out[2641]
  PIN rd_out[2642]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.405 0.070 874.475 ;
    END
  END rd_out[2642]
  PIN rd_out[2643]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.545 0.070 874.615 ;
    END
  END rd_out[2643]
  PIN rd_out[2644]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.685 0.070 874.755 ;
    END
  END rd_out[2644]
  PIN rd_out[2645]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.825 0.070 874.895 ;
    END
  END rd_out[2645]
  PIN rd_out[2646]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 874.965 0.070 875.035 ;
    END
  END rd_out[2646]
  PIN rd_out[2647]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.105 0.070 875.175 ;
    END
  END rd_out[2647]
  PIN rd_out[2648]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.245 0.070 875.315 ;
    END
  END rd_out[2648]
  PIN rd_out[2649]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.385 0.070 875.455 ;
    END
  END rd_out[2649]
  PIN rd_out[2650]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.525 0.070 875.595 ;
    END
  END rd_out[2650]
  PIN rd_out[2651]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.665 0.070 875.735 ;
    END
  END rd_out[2651]
  PIN rd_out[2652]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.805 0.070 875.875 ;
    END
  END rd_out[2652]
  PIN rd_out[2653]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 875.945 0.070 876.015 ;
    END
  END rd_out[2653]
  PIN rd_out[2654]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.085 0.070 876.155 ;
    END
  END rd_out[2654]
  PIN rd_out[2655]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.225 0.070 876.295 ;
    END
  END rd_out[2655]
  PIN rd_out[2656]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.365 0.070 876.435 ;
    END
  END rd_out[2656]
  PIN rd_out[2657]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.505 0.070 876.575 ;
    END
  END rd_out[2657]
  PIN rd_out[2658]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.645 0.070 876.715 ;
    END
  END rd_out[2658]
  PIN rd_out[2659]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.785 0.070 876.855 ;
    END
  END rd_out[2659]
  PIN rd_out[2660]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 876.925 0.070 876.995 ;
    END
  END rd_out[2660]
  PIN rd_out[2661]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.065 0.070 877.135 ;
    END
  END rd_out[2661]
  PIN rd_out[2662]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.205 0.070 877.275 ;
    END
  END rd_out[2662]
  PIN rd_out[2663]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.345 0.070 877.415 ;
    END
  END rd_out[2663]
  PIN rd_out[2664]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.485 0.070 877.555 ;
    END
  END rd_out[2664]
  PIN rd_out[2665]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.625 0.070 877.695 ;
    END
  END rd_out[2665]
  PIN rd_out[2666]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.765 0.070 877.835 ;
    END
  END rd_out[2666]
  PIN rd_out[2667]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 877.905 0.070 877.975 ;
    END
  END rd_out[2667]
  PIN rd_out[2668]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.045 0.070 878.115 ;
    END
  END rd_out[2668]
  PIN rd_out[2669]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.185 0.070 878.255 ;
    END
  END rd_out[2669]
  PIN rd_out[2670]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.325 0.070 878.395 ;
    END
  END rd_out[2670]
  PIN rd_out[2671]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.465 0.070 878.535 ;
    END
  END rd_out[2671]
  PIN rd_out[2672]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.605 0.070 878.675 ;
    END
  END rd_out[2672]
  PIN rd_out[2673]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.745 0.070 878.815 ;
    END
  END rd_out[2673]
  PIN rd_out[2674]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 878.885 0.070 878.955 ;
    END
  END rd_out[2674]
  PIN rd_out[2675]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.025 0.070 879.095 ;
    END
  END rd_out[2675]
  PIN rd_out[2676]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.165 0.070 879.235 ;
    END
  END rd_out[2676]
  PIN rd_out[2677]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.305 0.070 879.375 ;
    END
  END rd_out[2677]
  PIN rd_out[2678]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.445 0.070 879.515 ;
    END
  END rd_out[2678]
  PIN rd_out[2679]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.585 0.070 879.655 ;
    END
  END rd_out[2679]
  PIN rd_out[2680]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.725 0.070 879.795 ;
    END
  END rd_out[2680]
  PIN rd_out[2681]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 879.865 0.070 879.935 ;
    END
  END rd_out[2681]
  PIN rd_out[2682]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.005 0.070 880.075 ;
    END
  END rd_out[2682]
  PIN rd_out[2683]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.145 0.070 880.215 ;
    END
  END rd_out[2683]
  PIN rd_out[2684]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.285 0.070 880.355 ;
    END
  END rd_out[2684]
  PIN rd_out[2685]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.425 0.070 880.495 ;
    END
  END rd_out[2685]
  PIN rd_out[2686]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.565 0.070 880.635 ;
    END
  END rd_out[2686]
  PIN rd_out[2687]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.705 0.070 880.775 ;
    END
  END rd_out[2687]
  PIN rd_out[2688]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.845 0.070 880.915 ;
    END
  END rd_out[2688]
  PIN rd_out[2689]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 880.985 0.070 881.055 ;
    END
  END rd_out[2689]
  PIN rd_out[2690]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.125 0.070 881.195 ;
    END
  END rd_out[2690]
  PIN rd_out[2691]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.265 0.070 881.335 ;
    END
  END rd_out[2691]
  PIN rd_out[2692]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.405 0.070 881.475 ;
    END
  END rd_out[2692]
  PIN rd_out[2693]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.545 0.070 881.615 ;
    END
  END rd_out[2693]
  PIN rd_out[2694]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.685 0.070 881.755 ;
    END
  END rd_out[2694]
  PIN rd_out[2695]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.825 0.070 881.895 ;
    END
  END rd_out[2695]
  PIN rd_out[2696]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 881.965 0.070 882.035 ;
    END
  END rd_out[2696]
  PIN rd_out[2697]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.105 0.070 882.175 ;
    END
  END rd_out[2697]
  PIN rd_out[2698]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.245 0.070 882.315 ;
    END
  END rd_out[2698]
  PIN rd_out[2699]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.385 0.070 882.455 ;
    END
  END rd_out[2699]
  PIN rd_out[2700]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.525 0.070 882.595 ;
    END
  END rd_out[2700]
  PIN rd_out[2701]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.665 0.070 882.735 ;
    END
  END rd_out[2701]
  PIN rd_out[2702]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.805 0.070 882.875 ;
    END
  END rd_out[2702]
  PIN rd_out[2703]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 882.945 0.070 883.015 ;
    END
  END rd_out[2703]
  PIN rd_out[2704]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.085 0.070 883.155 ;
    END
  END rd_out[2704]
  PIN rd_out[2705]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.225 0.070 883.295 ;
    END
  END rd_out[2705]
  PIN rd_out[2706]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.365 0.070 883.435 ;
    END
  END rd_out[2706]
  PIN rd_out[2707]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.505 0.070 883.575 ;
    END
  END rd_out[2707]
  PIN rd_out[2708]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.645 0.070 883.715 ;
    END
  END rd_out[2708]
  PIN rd_out[2709]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.785 0.070 883.855 ;
    END
  END rd_out[2709]
  PIN rd_out[2710]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 883.925 0.070 883.995 ;
    END
  END rd_out[2710]
  PIN rd_out[2711]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.065 0.070 884.135 ;
    END
  END rd_out[2711]
  PIN rd_out[2712]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.205 0.070 884.275 ;
    END
  END rd_out[2712]
  PIN rd_out[2713]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.345 0.070 884.415 ;
    END
  END rd_out[2713]
  PIN rd_out[2714]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.485 0.070 884.555 ;
    END
  END rd_out[2714]
  PIN rd_out[2715]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.625 0.070 884.695 ;
    END
  END rd_out[2715]
  PIN rd_out[2716]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.765 0.070 884.835 ;
    END
  END rd_out[2716]
  PIN rd_out[2717]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 884.905 0.070 884.975 ;
    END
  END rd_out[2717]
  PIN rd_out[2718]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.045 0.070 885.115 ;
    END
  END rd_out[2718]
  PIN rd_out[2719]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.185 0.070 885.255 ;
    END
  END rd_out[2719]
  PIN rd_out[2720]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.325 0.070 885.395 ;
    END
  END rd_out[2720]
  PIN rd_out[2721]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.465 0.070 885.535 ;
    END
  END rd_out[2721]
  PIN rd_out[2722]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.605 0.070 885.675 ;
    END
  END rd_out[2722]
  PIN rd_out[2723]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.745 0.070 885.815 ;
    END
  END rd_out[2723]
  PIN rd_out[2724]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 885.885 0.070 885.955 ;
    END
  END rd_out[2724]
  PIN rd_out[2725]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.025 0.070 886.095 ;
    END
  END rd_out[2725]
  PIN rd_out[2726]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.165 0.070 886.235 ;
    END
  END rd_out[2726]
  PIN rd_out[2727]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.305 0.070 886.375 ;
    END
  END rd_out[2727]
  PIN rd_out[2728]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.445 0.070 886.515 ;
    END
  END rd_out[2728]
  PIN rd_out[2729]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.585 0.070 886.655 ;
    END
  END rd_out[2729]
  PIN rd_out[2730]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.725 0.070 886.795 ;
    END
  END rd_out[2730]
  PIN rd_out[2731]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 886.865 0.070 886.935 ;
    END
  END rd_out[2731]
  PIN rd_out[2732]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.005 0.070 887.075 ;
    END
  END rd_out[2732]
  PIN rd_out[2733]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.145 0.070 887.215 ;
    END
  END rd_out[2733]
  PIN rd_out[2734]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.285 0.070 887.355 ;
    END
  END rd_out[2734]
  PIN rd_out[2735]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.425 0.070 887.495 ;
    END
  END rd_out[2735]
  PIN rd_out[2736]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.565 0.070 887.635 ;
    END
  END rd_out[2736]
  PIN rd_out[2737]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.705 0.070 887.775 ;
    END
  END rd_out[2737]
  PIN rd_out[2738]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.845 0.070 887.915 ;
    END
  END rd_out[2738]
  PIN rd_out[2739]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 887.985 0.070 888.055 ;
    END
  END rd_out[2739]
  PIN rd_out[2740]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.125 0.070 888.195 ;
    END
  END rd_out[2740]
  PIN rd_out[2741]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.265 0.070 888.335 ;
    END
  END rd_out[2741]
  PIN rd_out[2742]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.405 0.070 888.475 ;
    END
  END rd_out[2742]
  PIN rd_out[2743]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.545 0.070 888.615 ;
    END
  END rd_out[2743]
  PIN rd_out[2744]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.685 0.070 888.755 ;
    END
  END rd_out[2744]
  PIN rd_out[2745]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.825 0.070 888.895 ;
    END
  END rd_out[2745]
  PIN rd_out[2746]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 888.965 0.070 889.035 ;
    END
  END rd_out[2746]
  PIN rd_out[2747]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.105 0.070 889.175 ;
    END
  END rd_out[2747]
  PIN rd_out[2748]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.245 0.070 889.315 ;
    END
  END rd_out[2748]
  PIN rd_out[2749]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.385 0.070 889.455 ;
    END
  END rd_out[2749]
  PIN rd_out[2750]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.525 0.070 889.595 ;
    END
  END rd_out[2750]
  PIN rd_out[2751]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.665 0.070 889.735 ;
    END
  END rd_out[2751]
  PIN rd_out[2752]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.805 0.070 889.875 ;
    END
  END rd_out[2752]
  PIN rd_out[2753]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 889.945 0.070 890.015 ;
    END
  END rd_out[2753]
  PIN rd_out[2754]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.085 0.070 890.155 ;
    END
  END rd_out[2754]
  PIN rd_out[2755]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.225 0.070 890.295 ;
    END
  END rd_out[2755]
  PIN rd_out[2756]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.365 0.070 890.435 ;
    END
  END rd_out[2756]
  PIN rd_out[2757]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.505 0.070 890.575 ;
    END
  END rd_out[2757]
  PIN rd_out[2758]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.645 0.070 890.715 ;
    END
  END rd_out[2758]
  PIN rd_out[2759]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.785 0.070 890.855 ;
    END
  END rd_out[2759]
  PIN rd_out[2760]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 890.925 0.070 890.995 ;
    END
  END rd_out[2760]
  PIN rd_out[2761]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.065 0.070 891.135 ;
    END
  END rd_out[2761]
  PIN rd_out[2762]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.205 0.070 891.275 ;
    END
  END rd_out[2762]
  PIN rd_out[2763]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.345 0.070 891.415 ;
    END
  END rd_out[2763]
  PIN rd_out[2764]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.485 0.070 891.555 ;
    END
  END rd_out[2764]
  PIN rd_out[2765]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.625 0.070 891.695 ;
    END
  END rd_out[2765]
  PIN rd_out[2766]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.765 0.070 891.835 ;
    END
  END rd_out[2766]
  PIN rd_out[2767]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 891.905 0.070 891.975 ;
    END
  END rd_out[2767]
  PIN rd_out[2768]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.045 0.070 892.115 ;
    END
  END rd_out[2768]
  PIN rd_out[2769]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.185 0.070 892.255 ;
    END
  END rd_out[2769]
  PIN rd_out[2770]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.325 0.070 892.395 ;
    END
  END rd_out[2770]
  PIN rd_out[2771]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.465 0.070 892.535 ;
    END
  END rd_out[2771]
  PIN rd_out[2772]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.605 0.070 892.675 ;
    END
  END rd_out[2772]
  PIN rd_out[2773]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.745 0.070 892.815 ;
    END
  END rd_out[2773]
  PIN rd_out[2774]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 892.885 0.070 892.955 ;
    END
  END rd_out[2774]
  PIN rd_out[2775]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.025 0.070 893.095 ;
    END
  END rd_out[2775]
  PIN rd_out[2776]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.165 0.070 893.235 ;
    END
  END rd_out[2776]
  PIN rd_out[2777]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.305 0.070 893.375 ;
    END
  END rd_out[2777]
  PIN rd_out[2778]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.445 0.070 893.515 ;
    END
  END rd_out[2778]
  PIN rd_out[2779]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.585 0.070 893.655 ;
    END
  END rd_out[2779]
  PIN rd_out[2780]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.725 0.070 893.795 ;
    END
  END rd_out[2780]
  PIN rd_out[2781]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 893.865 0.070 893.935 ;
    END
  END rd_out[2781]
  PIN rd_out[2782]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.005 0.070 894.075 ;
    END
  END rd_out[2782]
  PIN rd_out[2783]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.145 0.070 894.215 ;
    END
  END rd_out[2783]
  PIN rd_out[2784]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.285 0.070 894.355 ;
    END
  END rd_out[2784]
  PIN rd_out[2785]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.425 0.070 894.495 ;
    END
  END rd_out[2785]
  PIN rd_out[2786]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.565 0.070 894.635 ;
    END
  END rd_out[2786]
  PIN rd_out[2787]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.705 0.070 894.775 ;
    END
  END rd_out[2787]
  PIN rd_out[2788]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.845 0.070 894.915 ;
    END
  END rd_out[2788]
  PIN rd_out[2789]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 894.985 0.070 895.055 ;
    END
  END rd_out[2789]
  PIN rd_out[2790]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.125 0.070 895.195 ;
    END
  END rd_out[2790]
  PIN rd_out[2791]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.265 0.070 895.335 ;
    END
  END rd_out[2791]
  PIN rd_out[2792]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.405 0.070 895.475 ;
    END
  END rd_out[2792]
  PIN rd_out[2793]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.545 0.070 895.615 ;
    END
  END rd_out[2793]
  PIN rd_out[2794]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.685 0.070 895.755 ;
    END
  END rd_out[2794]
  PIN rd_out[2795]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.825 0.070 895.895 ;
    END
  END rd_out[2795]
  PIN rd_out[2796]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 895.965 0.070 896.035 ;
    END
  END rd_out[2796]
  PIN rd_out[2797]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.105 0.070 896.175 ;
    END
  END rd_out[2797]
  PIN rd_out[2798]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.245 0.070 896.315 ;
    END
  END rd_out[2798]
  PIN rd_out[2799]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.385 0.070 896.455 ;
    END
  END rd_out[2799]
  PIN rd_out[2800]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.525 0.070 896.595 ;
    END
  END rd_out[2800]
  PIN rd_out[2801]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.665 0.070 896.735 ;
    END
  END rd_out[2801]
  PIN rd_out[2802]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.805 0.070 896.875 ;
    END
  END rd_out[2802]
  PIN rd_out[2803]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 896.945 0.070 897.015 ;
    END
  END rd_out[2803]
  PIN rd_out[2804]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.085 0.070 897.155 ;
    END
  END rd_out[2804]
  PIN rd_out[2805]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.225 0.070 897.295 ;
    END
  END rd_out[2805]
  PIN rd_out[2806]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.365 0.070 897.435 ;
    END
  END rd_out[2806]
  PIN rd_out[2807]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.505 0.070 897.575 ;
    END
  END rd_out[2807]
  PIN rd_out[2808]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.645 0.070 897.715 ;
    END
  END rd_out[2808]
  PIN rd_out[2809]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.785 0.070 897.855 ;
    END
  END rd_out[2809]
  PIN rd_out[2810]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 897.925 0.070 897.995 ;
    END
  END rd_out[2810]
  PIN rd_out[2811]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.065 0.070 898.135 ;
    END
  END rd_out[2811]
  PIN rd_out[2812]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.205 0.070 898.275 ;
    END
  END rd_out[2812]
  PIN rd_out[2813]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.345 0.070 898.415 ;
    END
  END rd_out[2813]
  PIN rd_out[2814]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.485 0.070 898.555 ;
    END
  END rd_out[2814]
  PIN rd_out[2815]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.625 0.070 898.695 ;
    END
  END rd_out[2815]
  PIN rd_out[2816]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.765 0.070 898.835 ;
    END
  END rd_out[2816]
  PIN rd_out[2817]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 898.905 0.070 898.975 ;
    END
  END rd_out[2817]
  PIN rd_out[2818]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.045 0.070 899.115 ;
    END
  END rd_out[2818]
  PIN rd_out[2819]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.185 0.070 899.255 ;
    END
  END rd_out[2819]
  PIN rd_out[2820]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.325 0.070 899.395 ;
    END
  END rd_out[2820]
  PIN rd_out[2821]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.465 0.070 899.535 ;
    END
  END rd_out[2821]
  PIN rd_out[2822]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.605 0.070 899.675 ;
    END
  END rd_out[2822]
  PIN rd_out[2823]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.745 0.070 899.815 ;
    END
  END rd_out[2823]
  PIN rd_out[2824]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 899.885 0.070 899.955 ;
    END
  END rd_out[2824]
  PIN rd_out[2825]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.025 0.070 900.095 ;
    END
  END rd_out[2825]
  PIN rd_out[2826]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.165 0.070 900.235 ;
    END
  END rd_out[2826]
  PIN rd_out[2827]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.305 0.070 900.375 ;
    END
  END rd_out[2827]
  PIN rd_out[2828]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.445 0.070 900.515 ;
    END
  END rd_out[2828]
  PIN rd_out[2829]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.585 0.070 900.655 ;
    END
  END rd_out[2829]
  PIN rd_out[2830]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.725 0.070 900.795 ;
    END
  END rd_out[2830]
  PIN rd_out[2831]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 900.865 0.070 900.935 ;
    END
  END rd_out[2831]
  PIN rd_out[2832]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.005 0.070 901.075 ;
    END
  END rd_out[2832]
  PIN rd_out[2833]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.145 0.070 901.215 ;
    END
  END rd_out[2833]
  PIN rd_out[2834]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.285 0.070 901.355 ;
    END
  END rd_out[2834]
  PIN rd_out[2835]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.425 0.070 901.495 ;
    END
  END rd_out[2835]
  PIN rd_out[2836]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.565 0.070 901.635 ;
    END
  END rd_out[2836]
  PIN rd_out[2837]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.705 0.070 901.775 ;
    END
  END rd_out[2837]
  PIN rd_out[2838]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.845 0.070 901.915 ;
    END
  END rd_out[2838]
  PIN rd_out[2839]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 901.985 0.070 902.055 ;
    END
  END rd_out[2839]
  PIN rd_out[2840]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.125 0.070 902.195 ;
    END
  END rd_out[2840]
  PIN rd_out[2841]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.265 0.070 902.335 ;
    END
  END rd_out[2841]
  PIN rd_out[2842]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.405 0.070 902.475 ;
    END
  END rd_out[2842]
  PIN rd_out[2843]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.545 0.070 902.615 ;
    END
  END rd_out[2843]
  PIN rd_out[2844]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.685 0.070 902.755 ;
    END
  END rd_out[2844]
  PIN rd_out[2845]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.825 0.070 902.895 ;
    END
  END rd_out[2845]
  PIN rd_out[2846]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 902.965 0.070 903.035 ;
    END
  END rd_out[2846]
  PIN rd_out[2847]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 903.105 0.070 903.175 ;
    END
  END rd_out[2847]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1007.685 0.070 1007.755 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1007.825 0.070 1007.895 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1007.965 0.070 1008.035 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.105 0.070 1008.175 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.245 0.070 1008.315 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.385 0.070 1008.455 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.525 0.070 1008.595 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.665 0.070 1008.735 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.805 0.070 1008.875 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1008.945 0.070 1009.015 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1009.085 0.070 1009.155 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1009.225 0.070 1009.295 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1009.365 0.070 1009.435 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1009.505 0.070 1009.575 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1009.645 0.070 1009.715 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1009.785 0.070 1009.855 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1009.925 0.070 1009.995 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.065 0.070 1010.135 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.205 0.070 1010.275 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.345 0.070 1010.415 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.485 0.070 1010.555 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.625 0.070 1010.695 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.765 0.070 1010.835 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1010.905 0.070 1010.975 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1011.045 0.070 1011.115 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1011.185 0.070 1011.255 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1011.325 0.070 1011.395 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1011.465 0.070 1011.535 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1011.605 0.070 1011.675 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1011.745 0.070 1011.815 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1011.885 0.070 1011.955 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1012.025 0.070 1012.095 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1012.165 0.070 1012.235 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1012.305 0.070 1012.375 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1012.445 0.070 1012.515 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1012.585 0.070 1012.655 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1012.725 0.070 1012.795 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1012.865 0.070 1012.935 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.005 0.070 1013.075 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.145 0.070 1013.215 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.285 0.070 1013.355 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.425 0.070 1013.495 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.565 0.070 1013.635 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.705 0.070 1013.775 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.845 0.070 1013.915 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1013.985 0.070 1014.055 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.125 0.070 1014.195 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.265 0.070 1014.335 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.405 0.070 1014.475 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.545 0.070 1014.615 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.685 0.070 1014.755 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.825 0.070 1014.895 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1014.965 0.070 1015.035 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.105 0.070 1015.175 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.245 0.070 1015.315 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.385 0.070 1015.455 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.525 0.070 1015.595 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.665 0.070 1015.735 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.805 0.070 1015.875 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1015.945 0.070 1016.015 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1016.085 0.070 1016.155 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1016.225 0.070 1016.295 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1016.365 0.070 1016.435 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1016.505 0.070 1016.575 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1016.645 0.070 1016.715 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1016.785 0.070 1016.855 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1016.925 0.070 1016.995 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.065 0.070 1017.135 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.205 0.070 1017.275 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.345 0.070 1017.415 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.485 0.070 1017.555 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.625 0.070 1017.695 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.765 0.070 1017.835 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1017.905 0.070 1017.975 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1018.045 0.070 1018.115 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1018.185 0.070 1018.255 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1018.325 0.070 1018.395 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1018.465 0.070 1018.535 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1018.605 0.070 1018.675 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1018.745 0.070 1018.815 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1018.885 0.070 1018.955 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1019.025 0.070 1019.095 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1019.165 0.070 1019.235 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1019.305 0.070 1019.375 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1019.445 0.070 1019.515 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1019.585 0.070 1019.655 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1019.725 0.070 1019.795 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1019.865 0.070 1019.935 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.005 0.070 1020.075 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.145 0.070 1020.215 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.285 0.070 1020.355 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.425 0.070 1020.495 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.565 0.070 1020.635 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.705 0.070 1020.775 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.845 0.070 1020.915 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1020.985 0.070 1021.055 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1021.125 0.070 1021.195 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1021.265 0.070 1021.335 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1021.405 0.070 1021.475 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1021.545 0.070 1021.615 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1021.685 0.070 1021.755 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1021.825 0.070 1021.895 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1021.965 0.070 1022.035 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.105 0.070 1022.175 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.245 0.070 1022.315 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.385 0.070 1022.455 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.525 0.070 1022.595 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.665 0.070 1022.735 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.805 0.070 1022.875 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1022.945 0.070 1023.015 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1023.085 0.070 1023.155 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1023.225 0.070 1023.295 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1023.365 0.070 1023.435 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1023.505 0.070 1023.575 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1023.645 0.070 1023.715 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1023.785 0.070 1023.855 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1023.925 0.070 1023.995 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.065 0.070 1024.135 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.205 0.070 1024.275 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.345 0.070 1024.415 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.485 0.070 1024.555 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.625 0.070 1024.695 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.765 0.070 1024.835 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1024.905 0.070 1024.975 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1025.045 0.070 1025.115 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1025.185 0.070 1025.255 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1025.325 0.070 1025.395 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1025.465 0.070 1025.535 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1025.605 0.070 1025.675 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1025.745 0.070 1025.815 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1025.885 0.070 1025.955 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1026.025 0.070 1026.095 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1026.165 0.070 1026.235 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1026.305 0.070 1026.375 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1026.445 0.070 1026.515 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1026.585 0.070 1026.655 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1026.725 0.070 1026.795 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1026.865 0.070 1026.935 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.005 0.070 1027.075 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.145 0.070 1027.215 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.285 0.070 1027.355 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.425 0.070 1027.495 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.565 0.070 1027.635 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.705 0.070 1027.775 ;
    END
  END wd_in[143]
  PIN wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.845 0.070 1027.915 ;
    END
  END wd_in[144]
  PIN wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1027.985 0.070 1028.055 ;
    END
  END wd_in[145]
  PIN wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1028.125 0.070 1028.195 ;
    END
  END wd_in[146]
  PIN wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1028.265 0.070 1028.335 ;
    END
  END wd_in[147]
  PIN wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1028.405 0.070 1028.475 ;
    END
  END wd_in[148]
  PIN wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1028.545 0.070 1028.615 ;
    END
  END wd_in[149]
  PIN wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1028.685 0.070 1028.755 ;
    END
  END wd_in[150]
  PIN wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1028.825 0.070 1028.895 ;
    END
  END wd_in[151]
  PIN wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1028.965 0.070 1029.035 ;
    END
  END wd_in[152]
  PIN wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.105 0.070 1029.175 ;
    END
  END wd_in[153]
  PIN wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.245 0.070 1029.315 ;
    END
  END wd_in[154]
  PIN wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.385 0.070 1029.455 ;
    END
  END wd_in[155]
  PIN wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.525 0.070 1029.595 ;
    END
  END wd_in[156]
  PIN wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.665 0.070 1029.735 ;
    END
  END wd_in[157]
  PIN wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.805 0.070 1029.875 ;
    END
  END wd_in[158]
  PIN wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1029.945 0.070 1030.015 ;
    END
  END wd_in[159]
  PIN wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1030.085 0.070 1030.155 ;
    END
  END wd_in[160]
  PIN wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1030.225 0.070 1030.295 ;
    END
  END wd_in[161]
  PIN wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1030.365 0.070 1030.435 ;
    END
  END wd_in[162]
  PIN wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1030.505 0.070 1030.575 ;
    END
  END wd_in[163]
  PIN wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1030.645 0.070 1030.715 ;
    END
  END wd_in[164]
  PIN wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1030.785 0.070 1030.855 ;
    END
  END wd_in[165]
  PIN wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1030.925 0.070 1030.995 ;
    END
  END wd_in[166]
  PIN wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.065 0.070 1031.135 ;
    END
  END wd_in[167]
  PIN wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.205 0.070 1031.275 ;
    END
  END wd_in[168]
  PIN wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.345 0.070 1031.415 ;
    END
  END wd_in[169]
  PIN wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.485 0.070 1031.555 ;
    END
  END wd_in[170]
  PIN wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.625 0.070 1031.695 ;
    END
  END wd_in[171]
  PIN wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.765 0.070 1031.835 ;
    END
  END wd_in[172]
  PIN wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1031.905 0.070 1031.975 ;
    END
  END wd_in[173]
  PIN wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1032.045 0.070 1032.115 ;
    END
  END wd_in[174]
  PIN wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1032.185 0.070 1032.255 ;
    END
  END wd_in[175]
  PIN wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1032.325 0.070 1032.395 ;
    END
  END wd_in[176]
  PIN wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1032.465 0.070 1032.535 ;
    END
  END wd_in[177]
  PIN wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1032.605 0.070 1032.675 ;
    END
  END wd_in[178]
  PIN wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1032.745 0.070 1032.815 ;
    END
  END wd_in[179]
  PIN wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1032.885 0.070 1032.955 ;
    END
  END wd_in[180]
  PIN wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1033.025 0.070 1033.095 ;
    END
  END wd_in[181]
  PIN wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1033.165 0.070 1033.235 ;
    END
  END wd_in[182]
  PIN wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1033.305 0.070 1033.375 ;
    END
  END wd_in[183]
  PIN wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1033.445 0.070 1033.515 ;
    END
  END wd_in[184]
  PIN wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1033.585 0.070 1033.655 ;
    END
  END wd_in[185]
  PIN wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1033.725 0.070 1033.795 ;
    END
  END wd_in[186]
  PIN wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1033.865 0.070 1033.935 ;
    END
  END wd_in[187]
  PIN wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.005 0.070 1034.075 ;
    END
  END wd_in[188]
  PIN wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.145 0.070 1034.215 ;
    END
  END wd_in[189]
  PIN wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.285 0.070 1034.355 ;
    END
  END wd_in[190]
  PIN wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.425 0.070 1034.495 ;
    END
  END wd_in[191]
  PIN wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.565 0.070 1034.635 ;
    END
  END wd_in[192]
  PIN wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.705 0.070 1034.775 ;
    END
  END wd_in[193]
  PIN wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.845 0.070 1034.915 ;
    END
  END wd_in[194]
  PIN wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1034.985 0.070 1035.055 ;
    END
  END wd_in[195]
  PIN wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.125 0.070 1035.195 ;
    END
  END wd_in[196]
  PIN wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.265 0.070 1035.335 ;
    END
  END wd_in[197]
  PIN wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.405 0.070 1035.475 ;
    END
  END wd_in[198]
  PIN wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.545 0.070 1035.615 ;
    END
  END wd_in[199]
  PIN wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.685 0.070 1035.755 ;
    END
  END wd_in[200]
  PIN wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.825 0.070 1035.895 ;
    END
  END wd_in[201]
  PIN wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1035.965 0.070 1036.035 ;
    END
  END wd_in[202]
  PIN wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.105 0.070 1036.175 ;
    END
  END wd_in[203]
  PIN wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.245 0.070 1036.315 ;
    END
  END wd_in[204]
  PIN wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.385 0.070 1036.455 ;
    END
  END wd_in[205]
  PIN wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.525 0.070 1036.595 ;
    END
  END wd_in[206]
  PIN wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.665 0.070 1036.735 ;
    END
  END wd_in[207]
  PIN wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.805 0.070 1036.875 ;
    END
  END wd_in[208]
  PIN wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1036.945 0.070 1037.015 ;
    END
  END wd_in[209]
  PIN wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1037.085 0.070 1037.155 ;
    END
  END wd_in[210]
  PIN wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1037.225 0.070 1037.295 ;
    END
  END wd_in[211]
  PIN wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1037.365 0.070 1037.435 ;
    END
  END wd_in[212]
  PIN wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1037.505 0.070 1037.575 ;
    END
  END wd_in[213]
  PIN wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1037.645 0.070 1037.715 ;
    END
  END wd_in[214]
  PIN wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1037.785 0.070 1037.855 ;
    END
  END wd_in[215]
  PIN wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1037.925 0.070 1037.995 ;
    END
  END wd_in[216]
  PIN wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.065 0.070 1038.135 ;
    END
  END wd_in[217]
  PIN wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.205 0.070 1038.275 ;
    END
  END wd_in[218]
  PIN wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.345 0.070 1038.415 ;
    END
  END wd_in[219]
  PIN wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.485 0.070 1038.555 ;
    END
  END wd_in[220]
  PIN wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.625 0.070 1038.695 ;
    END
  END wd_in[221]
  PIN wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.765 0.070 1038.835 ;
    END
  END wd_in[222]
  PIN wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1038.905 0.070 1038.975 ;
    END
  END wd_in[223]
  PIN wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1039.045 0.070 1039.115 ;
    END
  END wd_in[224]
  PIN wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1039.185 0.070 1039.255 ;
    END
  END wd_in[225]
  PIN wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1039.325 0.070 1039.395 ;
    END
  END wd_in[226]
  PIN wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1039.465 0.070 1039.535 ;
    END
  END wd_in[227]
  PIN wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1039.605 0.070 1039.675 ;
    END
  END wd_in[228]
  PIN wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1039.745 0.070 1039.815 ;
    END
  END wd_in[229]
  PIN wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1039.885 0.070 1039.955 ;
    END
  END wd_in[230]
  PIN wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1040.025 0.070 1040.095 ;
    END
  END wd_in[231]
  PIN wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1040.165 0.070 1040.235 ;
    END
  END wd_in[232]
  PIN wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1040.305 0.070 1040.375 ;
    END
  END wd_in[233]
  PIN wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1040.445 0.070 1040.515 ;
    END
  END wd_in[234]
  PIN wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1040.585 0.070 1040.655 ;
    END
  END wd_in[235]
  PIN wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1040.725 0.070 1040.795 ;
    END
  END wd_in[236]
  PIN wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1040.865 0.070 1040.935 ;
    END
  END wd_in[237]
  PIN wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.005 0.070 1041.075 ;
    END
  END wd_in[238]
  PIN wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.145 0.070 1041.215 ;
    END
  END wd_in[239]
  PIN wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.285 0.070 1041.355 ;
    END
  END wd_in[240]
  PIN wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.425 0.070 1041.495 ;
    END
  END wd_in[241]
  PIN wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.565 0.070 1041.635 ;
    END
  END wd_in[242]
  PIN wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.705 0.070 1041.775 ;
    END
  END wd_in[243]
  PIN wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.845 0.070 1041.915 ;
    END
  END wd_in[244]
  PIN wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1041.985 0.070 1042.055 ;
    END
  END wd_in[245]
  PIN wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1042.125 0.070 1042.195 ;
    END
  END wd_in[246]
  PIN wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1042.265 0.070 1042.335 ;
    END
  END wd_in[247]
  PIN wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1042.405 0.070 1042.475 ;
    END
  END wd_in[248]
  PIN wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1042.545 0.070 1042.615 ;
    END
  END wd_in[249]
  PIN wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1042.685 0.070 1042.755 ;
    END
  END wd_in[250]
  PIN wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1042.825 0.070 1042.895 ;
    END
  END wd_in[251]
  PIN wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1042.965 0.070 1043.035 ;
    END
  END wd_in[252]
  PIN wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.105 0.070 1043.175 ;
    END
  END wd_in[253]
  PIN wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.245 0.070 1043.315 ;
    END
  END wd_in[254]
  PIN wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.385 0.070 1043.455 ;
    END
  END wd_in[255]
  PIN wd_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.525 0.070 1043.595 ;
    END
  END wd_in[256]
  PIN wd_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.665 0.070 1043.735 ;
    END
  END wd_in[257]
  PIN wd_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.805 0.070 1043.875 ;
    END
  END wd_in[258]
  PIN wd_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1043.945 0.070 1044.015 ;
    END
  END wd_in[259]
  PIN wd_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1044.085 0.070 1044.155 ;
    END
  END wd_in[260]
  PIN wd_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1044.225 0.070 1044.295 ;
    END
  END wd_in[261]
  PIN wd_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1044.365 0.070 1044.435 ;
    END
  END wd_in[262]
  PIN wd_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1044.505 0.070 1044.575 ;
    END
  END wd_in[263]
  PIN wd_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1044.645 0.070 1044.715 ;
    END
  END wd_in[264]
  PIN wd_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1044.785 0.070 1044.855 ;
    END
  END wd_in[265]
  PIN wd_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1044.925 0.070 1044.995 ;
    END
  END wd_in[266]
  PIN wd_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.065 0.070 1045.135 ;
    END
  END wd_in[267]
  PIN wd_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.205 0.070 1045.275 ;
    END
  END wd_in[268]
  PIN wd_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.345 0.070 1045.415 ;
    END
  END wd_in[269]
  PIN wd_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.485 0.070 1045.555 ;
    END
  END wd_in[270]
  PIN wd_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.625 0.070 1045.695 ;
    END
  END wd_in[271]
  PIN wd_in[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.765 0.070 1045.835 ;
    END
  END wd_in[272]
  PIN wd_in[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1045.905 0.070 1045.975 ;
    END
  END wd_in[273]
  PIN wd_in[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.045 0.070 1046.115 ;
    END
  END wd_in[274]
  PIN wd_in[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.185 0.070 1046.255 ;
    END
  END wd_in[275]
  PIN wd_in[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.325 0.070 1046.395 ;
    END
  END wd_in[276]
  PIN wd_in[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.465 0.070 1046.535 ;
    END
  END wd_in[277]
  PIN wd_in[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.605 0.070 1046.675 ;
    END
  END wd_in[278]
  PIN wd_in[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.745 0.070 1046.815 ;
    END
  END wd_in[279]
  PIN wd_in[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1046.885 0.070 1046.955 ;
    END
  END wd_in[280]
  PIN wd_in[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1047.025 0.070 1047.095 ;
    END
  END wd_in[281]
  PIN wd_in[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1047.165 0.070 1047.235 ;
    END
  END wd_in[282]
  PIN wd_in[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1047.305 0.070 1047.375 ;
    END
  END wd_in[283]
  PIN wd_in[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1047.445 0.070 1047.515 ;
    END
  END wd_in[284]
  PIN wd_in[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1047.585 0.070 1047.655 ;
    END
  END wd_in[285]
  PIN wd_in[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1047.725 0.070 1047.795 ;
    END
  END wd_in[286]
  PIN wd_in[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1047.865 0.070 1047.935 ;
    END
  END wd_in[287]
  PIN wd_in[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.005 0.070 1048.075 ;
    END
  END wd_in[288]
  PIN wd_in[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.145 0.070 1048.215 ;
    END
  END wd_in[289]
  PIN wd_in[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.285 0.070 1048.355 ;
    END
  END wd_in[290]
  PIN wd_in[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.425 0.070 1048.495 ;
    END
  END wd_in[291]
  PIN wd_in[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.565 0.070 1048.635 ;
    END
  END wd_in[292]
  PIN wd_in[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.705 0.070 1048.775 ;
    END
  END wd_in[293]
  PIN wd_in[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.845 0.070 1048.915 ;
    END
  END wd_in[294]
  PIN wd_in[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1048.985 0.070 1049.055 ;
    END
  END wd_in[295]
  PIN wd_in[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1049.125 0.070 1049.195 ;
    END
  END wd_in[296]
  PIN wd_in[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1049.265 0.070 1049.335 ;
    END
  END wd_in[297]
  PIN wd_in[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1049.405 0.070 1049.475 ;
    END
  END wd_in[298]
  PIN wd_in[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1049.545 0.070 1049.615 ;
    END
  END wd_in[299]
  PIN wd_in[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1049.685 0.070 1049.755 ;
    END
  END wd_in[300]
  PIN wd_in[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1049.825 0.070 1049.895 ;
    END
  END wd_in[301]
  PIN wd_in[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1049.965 0.070 1050.035 ;
    END
  END wd_in[302]
  PIN wd_in[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.105 0.070 1050.175 ;
    END
  END wd_in[303]
  PIN wd_in[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.245 0.070 1050.315 ;
    END
  END wd_in[304]
  PIN wd_in[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.385 0.070 1050.455 ;
    END
  END wd_in[305]
  PIN wd_in[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.525 0.070 1050.595 ;
    END
  END wd_in[306]
  PIN wd_in[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.665 0.070 1050.735 ;
    END
  END wd_in[307]
  PIN wd_in[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.805 0.070 1050.875 ;
    END
  END wd_in[308]
  PIN wd_in[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1050.945 0.070 1051.015 ;
    END
  END wd_in[309]
  PIN wd_in[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1051.085 0.070 1051.155 ;
    END
  END wd_in[310]
  PIN wd_in[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1051.225 0.070 1051.295 ;
    END
  END wd_in[311]
  PIN wd_in[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1051.365 0.070 1051.435 ;
    END
  END wd_in[312]
  PIN wd_in[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1051.505 0.070 1051.575 ;
    END
  END wd_in[313]
  PIN wd_in[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1051.645 0.070 1051.715 ;
    END
  END wd_in[314]
  PIN wd_in[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1051.785 0.070 1051.855 ;
    END
  END wd_in[315]
  PIN wd_in[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1051.925 0.070 1051.995 ;
    END
  END wd_in[316]
  PIN wd_in[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.065 0.070 1052.135 ;
    END
  END wd_in[317]
  PIN wd_in[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.205 0.070 1052.275 ;
    END
  END wd_in[318]
  PIN wd_in[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.345 0.070 1052.415 ;
    END
  END wd_in[319]
  PIN wd_in[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.485 0.070 1052.555 ;
    END
  END wd_in[320]
  PIN wd_in[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.625 0.070 1052.695 ;
    END
  END wd_in[321]
  PIN wd_in[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.765 0.070 1052.835 ;
    END
  END wd_in[322]
  PIN wd_in[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1052.905 0.070 1052.975 ;
    END
  END wd_in[323]
  PIN wd_in[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1053.045 0.070 1053.115 ;
    END
  END wd_in[324]
  PIN wd_in[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1053.185 0.070 1053.255 ;
    END
  END wd_in[325]
  PIN wd_in[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1053.325 0.070 1053.395 ;
    END
  END wd_in[326]
  PIN wd_in[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1053.465 0.070 1053.535 ;
    END
  END wd_in[327]
  PIN wd_in[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1053.605 0.070 1053.675 ;
    END
  END wd_in[328]
  PIN wd_in[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1053.745 0.070 1053.815 ;
    END
  END wd_in[329]
  PIN wd_in[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1053.885 0.070 1053.955 ;
    END
  END wd_in[330]
  PIN wd_in[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1054.025 0.070 1054.095 ;
    END
  END wd_in[331]
  PIN wd_in[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1054.165 0.070 1054.235 ;
    END
  END wd_in[332]
  PIN wd_in[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1054.305 0.070 1054.375 ;
    END
  END wd_in[333]
  PIN wd_in[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1054.445 0.070 1054.515 ;
    END
  END wd_in[334]
  PIN wd_in[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1054.585 0.070 1054.655 ;
    END
  END wd_in[335]
  PIN wd_in[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1054.725 0.070 1054.795 ;
    END
  END wd_in[336]
  PIN wd_in[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1054.865 0.070 1054.935 ;
    END
  END wd_in[337]
  PIN wd_in[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.005 0.070 1055.075 ;
    END
  END wd_in[338]
  PIN wd_in[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.145 0.070 1055.215 ;
    END
  END wd_in[339]
  PIN wd_in[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.285 0.070 1055.355 ;
    END
  END wd_in[340]
  PIN wd_in[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.425 0.070 1055.495 ;
    END
  END wd_in[341]
  PIN wd_in[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.565 0.070 1055.635 ;
    END
  END wd_in[342]
  PIN wd_in[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.705 0.070 1055.775 ;
    END
  END wd_in[343]
  PIN wd_in[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.845 0.070 1055.915 ;
    END
  END wd_in[344]
  PIN wd_in[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1055.985 0.070 1056.055 ;
    END
  END wd_in[345]
  PIN wd_in[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1056.125 0.070 1056.195 ;
    END
  END wd_in[346]
  PIN wd_in[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1056.265 0.070 1056.335 ;
    END
  END wd_in[347]
  PIN wd_in[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1056.405 0.070 1056.475 ;
    END
  END wd_in[348]
  PIN wd_in[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1056.545 0.070 1056.615 ;
    END
  END wd_in[349]
  PIN wd_in[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1056.685 0.070 1056.755 ;
    END
  END wd_in[350]
  PIN wd_in[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1056.825 0.070 1056.895 ;
    END
  END wd_in[351]
  PIN wd_in[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1056.965 0.070 1057.035 ;
    END
  END wd_in[352]
  PIN wd_in[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.105 0.070 1057.175 ;
    END
  END wd_in[353]
  PIN wd_in[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.245 0.070 1057.315 ;
    END
  END wd_in[354]
  PIN wd_in[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.385 0.070 1057.455 ;
    END
  END wd_in[355]
  PIN wd_in[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.525 0.070 1057.595 ;
    END
  END wd_in[356]
  PIN wd_in[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.665 0.070 1057.735 ;
    END
  END wd_in[357]
  PIN wd_in[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.805 0.070 1057.875 ;
    END
  END wd_in[358]
  PIN wd_in[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1057.945 0.070 1058.015 ;
    END
  END wd_in[359]
  PIN wd_in[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1058.085 0.070 1058.155 ;
    END
  END wd_in[360]
  PIN wd_in[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1058.225 0.070 1058.295 ;
    END
  END wd_in[361]
  PIN wd_in[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1058.365 0.070 1058.435 ;
    END
  END wd_in[362]
  PIN wd_in[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1058.505 0.070 1058.575 ;
    END
  END wd_in[363]
  PIN wd_in[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1058.645 0.070 1058.715 ;
    END
  END wd_in[364]
  PIN wd_in[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1058.785 0.070 1058.855 ;
    END
  END wd_in[365]
  PIN wd_in[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1058.925 0.070 1058.995 ;
    END
  END wd_in[366]
  PIN wd_in[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.065 0.070 1059.135 ;
    END
  END wd_in[367]
  PIN wd_in[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.205 0.070 1059.275 ;
    END
  END wd_in[368]
  PIN wd_in[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.345 0.070 1059.415 ;
    END
  END wd_in[369]
  PIN wd_in[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.485 0.070 1059.555 ;
    END
  END wd_in[370]
  PIN wd_in[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.625 0.070 1059.695 ;
    END
  END wd_in[371]
  PIN wd_in[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.765 0.070 1059.835 ;
    END
  END wd_in[372]
  PIN wd_in[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1059.905 0.070 1059.975 ;
    END
  END wd_in[373]
  PIN wd_in[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1060.045 0.070 1060.115 ;
    END
  END wd_in[374]
  PIN wd_in[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1060.185 0.070 1060.255 ;
    END
  END wd_in[375]
  PIN wd_in[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1060.325 0.070 1060.395 ;
    END
  END wd_in[376]
  PIN wd_in[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1060.465 0.070 1060.535 ;
    END
  END wd_in[377]
  PIN wd_in[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1060.605 0.070 1060.675 ;
    END
  END wd_in[378]
  PIN wd_in[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1060.745 0.070 1060.815 ;
    END
  END wd_in[379]
  PIN wd_in[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1060.885 0.070 1060.955 ;
    END
  END wd_in[380]
  PIN wd_in[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1061.025 0.070 1061.095 ;
    END
  END wd_in[381]
  PIN wd_in[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1061.165 0.070 1061.235 ;
    END
  END wd_in[382]
  PIN wd_in[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1061.305 0.070 1061.375 ;
    END
  END wd_in[383]
  PIN wd_in[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1061.445 0.070 1061.515 ;
    END
  END wd_in[384]
  PIN wd_in[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1061.585 0.070 1061.655 ;
    END
  END wd_in[385]
  PIN wd_in[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1061.725 0.070 1061.795 ;
    END
  END wd_in[386]
  PIN wd_in[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1061.865 0.070 1061.935 ;
    END
  END wd_in[387]
  PIN wd_in[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.005 0.070 1062.075 ;
    END
  END wd_in[388]
  PIN wd_in[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.145 0.070 1062.215 ;
    END
  END wd_in[389]
  PIN wd_in[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.285 0.070 1062.355 ;
    END
  END wd_in[390]
  PIN wd_in[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.425 0.070 1062.495 ;
    END
  END wd_in[391]
  PIN wd_in[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.565 0.070 1062.635 ;
    END
  END wd_in[392]
  PIN wd_in[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.705 0.070 1062.775 ;
    END
  END wd_in[393]
  PIN wd_in[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.845 0.070 1062.915 ;
    END
  END wd_in[394]
  PIN wd_in[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1062.985 0.070 1063.055 ;
    END
  END wd_in[395]
  PIN wd_in[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1063.125 0.070 1063.195 ;
    END
  END wd_in[396]
  PIN wd_in[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1063.265 0.070 1063.335 ;
    END
  END wd_in[397]
  PIN wd_in[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1063.405 0.070 1063.475 ;
    END
  END wd_in[398]
  PIN wd_in[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1063.545 0.070 1063.615 ;
    END
  END wd_in[399]
  PIN wd_in[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1063.685 0.070 1063.755 ;
    END
  END wd_in[400]
  PIN wd_in[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1063.825 0.070 1063.895 ;
    END
  END wd_in[401]
  PIN wd_in[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1063.965 0.070 1064.035 ;
    END
  END wd_in[402]
  PIN wd_in[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.105 0.070 1064.175 ;
    END
  END wd_in[403]
  PIN wd_in[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.245 0.070 1064.315 ;
    END
  END wd_in[404]
  PIN wd_in[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.385 0.070 1064.455 ;
    END
  END wd_in[405]
  PIN wd_in[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.525 0.070 1064.595 ;
    END
  END wd_in[406]
  PIN wd_in[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.665 0.070 1064.735 ;
    END
  END wd_in[407]
  PIN wd_in[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.805 0.070 1064.875 ;
    END
  END wd_in[408]
  PIN wd_in[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1064.945 0.070 1065.015 ;
    END
  END wd_in[409]
  PIN wd_in[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1065.085 0.070 1065.155 ;
    END
  END wd_in[410]
  PIN wd_in[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1065.225 0.070 1065.295 ;
    END
  END wd_in[411]
  PIN wd_in[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1065.365 0.070 1065.435 ;
    END
  END wd_in[412]
  PIN wd_in[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1065.505 0.070 1065.575 ;
    END
  END wd_in[413]
  PIN wd_in[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1065.645 0.070 1065.715 ;
    END
  END wd_in[414]
  PIN wd_in[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1065.785 0.070 1065.855 ;
    END
  END wd_in[415]
  PIN wd_in[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1065.925 0.070 1065.995 ;
    END
  END wd_in[416]
  PIN wd_in[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.065 0.070 1066.135 ;
    END
  END wd_in[417]
  PIN wd_in[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.205 0.070 1066.275 ;
    END
  END wd_in[418]
  PIN wd_in[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.345 0.070 1066.415 ;
    END
  END wd_in[419]
  PIN wd_in[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.485 0.070 1066.555 ;
    END
  END wd_in[420]
  PIN wd_in[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.625 0.070 1066.695 ;
    END
  END wd_in[421]
  PIN wd_in[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.765 0.070 1066.835 ;
    END
  END wd_in[422]
  PIN wd_in[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1066.905 0.070 1066.975 ;
    END
  END wd_in[423]
  PIN wd_in[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1067.045 0.070 1067.115 ;
    END
  END wd_in[424]
  PIN wd_in[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1067.185 0.070 1067.255 ;
    END
  END wd_in[425]
  PIN wd_in[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1067.325 0.070 1067.395 ;
    END
  END wd_in[426]
  PIN wd_in[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1067.465 0.070 1067.535 ;
    END
  END wd_in[427]
  PIN wd_in[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1067.605 0.070 1067.675 ;
    END
  END wd_in[428]
  PIN wd_in[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1067.745 0.070 1067.815 ;
    END
  END wd_in[429]
  PIN wd_in[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1067.885 0.070 1067.955 ;
    END
  END wd_in[430]
  PIN wd_in[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.025 0.070 1068.095 ;
    END
  END wd_in[431]
  PIN wd_in[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.165 0.070 1068.235 ;
    END
  END wd_in[432]
  PIN wd_in[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.305 0.070 1068.375 ;
    END
  END wd_in[433]
  PIN wd_in[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.445 0.070 1068.515 ;
    END
  END wd_in[434]
  PIN wd_in[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.585 0.070 1068.655 ;
    END
  END wd_in[435]
  PIN wd_in[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.725 0.070 1068.795 ;
    END
  END wd_in[436]
  PIN wd_in[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1068.865 0.070 1068.935 ;
    END
  END wd_in[437]
  PIN wd_in[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.005 0.070 1069.075 ;
    END
  END wd_in[438]
  PIN wd_in[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.145 0.070 1069.215 ;
    END
  END wd_in[439]
  PIN wd_in[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.285 0.070 1069.355 ;
    END
  END wd_in[440]
  PIN wd_in[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.425 0.070 1069.495 ;
    END
  END wd_in[441]
  PIN wd_in[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.565 0.070 1069.635 ;
    END
  END wd_in[442]
  PIN wd_in[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.705 0.070 1069.775 ;
    END
  END wd_in[443]
  PIN wd_in[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.845 0.070 1069.915 ;
    END
  END wd_in[444]
  PIN wd_in[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1069.985 0.070 1070.055 ;
    END
  END wd_in[445]
  PIN wd_in[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1070.125 0.070 1070.195 ;
    END
  END wd_in[446]
  PIN wd_in[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1070.265 0.070 1070.335 ;
    END
  END wd_in[447]
  PIN wd_in[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1070.405 0.070 1070.475 ;
    END
  END wd_in[448]
  PIN wd_in[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1070.545 0.070 1070.615 ;
    END
  END wd_in[449]
  PIN wd_in[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1070.685 0.070 1070.755 ;
    END
  END wd_in[450]
  PIN wd_in[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1070.825 0.070 1070.895 ;
    END
  END wd_in[451]
  PIN wd_in[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1070.965 0.070 1071.035 ;
    END
  END wd_in[452]
  PIN wd_in[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.105 0.070 1071.175 ;
    END
  END wd_in[453]
  PIN wd_in[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.245 0.070 1071.315 ;
    END
  END wd_in[454]
  PIN wd_in[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.385 0.070 1071.455 ;
    END
  END wd_in[455]
  PIN wd_in[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.525 0.070 1071.595 ;
    END
  END wd_in[456]
  PIN wd_in[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.665 0.070 1071.735 ;
    END
  END wd_in[457]
  PIN wd_in[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.805 0.070 1071.875 ;
    END
  END wd_in[458]
  PIN wd_in[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1071.945 0.070 1072.015 ;
    END
  END wd_in[459]
  PIN wd_in[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1072.085 0.070 1072.155 ;
    END
  END wd_in[460]
  PIN wd_in[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1072.225 0.070 1072.295 ;
    END
  END wd_in[461]
  PIN wd_in[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1072.365 0.070 1072.435 ;
    END
  END wd_in[462]
  PIN wd_in[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1072.505 0.070 1072.575 ;
    END
  END wd_in[463]
  PIN wd_in[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1072.645 0.070 1072.715 ;
    END
  END wd_in[464]
  PIN wd_in[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1072.785 0.070 1072.855 ;
    END
  END wd_in[465]
  PIN wd_in[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1072.925 0.070 1072.995 ;
    END
  END wd_in[466]
  PIN wd_in[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.065 0.070 1073.135 ;
    END
  END wd_in[467]
  PIN wd_in[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.205 0.070 1073.275 ;
    END
  END wd_in[468]
  PIN wd_in[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.345 0.070 1073.415 ;
    END
  END wd_in[469]
  PIN wd_in[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.485 0.070 1073.555 ;
    END
  END wd_in[470]
  PIN wd_in[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.625 0.070 1073.695 ;
    END
  END wd_in[471]
  PIN wd_in[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.765 0.070 1073.835 ;
    END
  END wd_in[472]
  PIN wd_in[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1073.905 0.070 1073.975 ;
    END
  END wd_in[473]
  PIN wd_in[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1074.045 0.070 1074.115 ;
    END
  END wd_in[474]
  PIN wd_in[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1074.185 0.070 1074.255 ;
    END
  END wd_in[475]
  PIN wd_in[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1074.325 0.070 1074.395 ;
    END
  END wd_in[476]
  PIN wd_in[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1074.465 0.070 1074.535 ;
    END
  END wd_in[477]
  PIN wd_in[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1074.605 0.070 1074.675 ;
    END
  END wd_in[478]
  PIN wd_in[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1074.745 0.070 1074.815 ;
    END
  END wd_in[479]
  PIN wd_in[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1074.885 0.070 1074.955 ;
    END
  END wd_in[480]
  PIN wd_in[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1075.025 0.070 1075.095 ;
    END
  END wd_in[481]
  PIN wd_in[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1075.165 0.070 1075.235 ;
    END
  END wd_in[482]
  PIN wd_in[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1075.305 0.070 1075.375 ;
    END
  END wd_in[483]
  PIN wd_in[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1075.445 0.070 1075.515 ;
    END
  END wd_in[484]
  PIN wd_in[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1075.585 0.070 1075.655 ;
    END
  END wd_in[485]
  PIN wd_in[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1075.725 0.070 1075.795 ;
    END
  END wd_in[486]
  PIN wd_in[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1075.865 0.070 1075.935 ;
    END
  END wd_in[487]
  PIN wd_in[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.005 0.070 1076.075 ;
    END
  END wd_in[488]
  PIN wd_in[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.145 0.070 1076.215 ;
    END
  END wd_in[489]
  PIN wd_in[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.285 0.070 1076.355 ;
    END
  END wd_in[490]
  PIN wd_in[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.425 0.070 1076.495 ;
    END
  END wd_in[491]
  PIN wd_in[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.565 0.070 1076.635 ;
    END
  END wd_in[492]
  PIN wd_in[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.705 0.070 1076.775 ;
    END
  END wd_in[493]
  PIN wd_in[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.845 0.070 1076.915 ;
    END
  END wd_in[494]
  PIN wd_in[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1076.985 0.070 1077.055 ;
    END
  END wd_in[495]
  PIN wd_in[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1077.125 0.070 1077.195 ;
    END
  END wd_in[496]
  PIN wd_in[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1077.265 0.070 1077.335 ;
    END
  END wd_in[497]
  PIN wd_in[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1077.405 0.070 1077.475 ;
    END
  END wd_in[498]
  PIN wd_in[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1077.545 0.070 1077.615 ;
    END
  END wd_in[499]
  PIN wd_in[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1077.685 0.070 1077.755 ;
    END
  END wd_in[500]
  PIN wd_in[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1077.825 0.070 1077.895 ;
    END
  END wd_in[501]
  PIN wd_in[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1077.965 0.070 1078.035 ;
    END
  END wd_in[502]
  PIN wd_in[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.105 0.070 1078.175 ;
    END
  END wd_in[503]
  PIN wd_in[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.245 0.070 1078.315 ;
    END
  END wd_in[504]
  PIN wd_in[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.385 0.070 1078.455 ;
    END
  END wd_in[505]
  PIN wd_in[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.525 0.070 1078.595 ;
    END
  END wd_in[506]
  PIN wd_in[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.665 0.070 1078.735 ;
    END
  END wd_in[507]
  PIN wd_in[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.805 0.070 1078.875 ;
    END
  END wd_in[508]
  PIN wd_in[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1078.945 0.070 1079.015 ;
    END
  END wd_in[509]
  PIN wd_in[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1079.085 0.070 1079.155 ;
    END
  END wd_in[510]
  PIN wd_in[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1079.225 0.070 1079.295 ;
    END
  END wd_in[511]
  PIN wd_in[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1079.365 0.070 1079.435 ;
    END
  END wd_in[512]
  PIN wd_in[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1079.505 0.070 1079.575 ;
    END
  END wd_in[513]
  PIN wd_in[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1079.645 0.070 1079.715 ;
    END
  END wd_in[514]
  PIN wd_in[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1079.785 0.070 1079.855 ;
    END
  END wd_in[515]
  PIN wd_in[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1079.925 0.070 1079.995 ;
    END
  END wd_in[516]
  PIN wd_in[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.065 0.070 1080.135 ;
    END
  END wd_in[517]
  PIN wd_in[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.205 0.070 1080.275 ;
    END
  END wd_in[518]
  PIN wd_in[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.345 0.070 1080.415 ;
    END
  END wd_in[519]
  PIN wd_in[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.485 0.070 1080.555 ;
    END
  END wd_in[520]
  PIN wd_in[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.625 0.070 1080.695 ;
    END
  END wd_in[521]
  PIN wd_in[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.765 0.070 1080.835 ;
    END
  END wd_in[522]
  PIN wd_in[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1080.905 0.070 1080.975 ;
    END
  END wd_in[523]
  PIN wd_in[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1081.045 0.070 1081.115 ;
    END
  END wd_in[524]
  PIN wd_in[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1081.185 0.070 1081.255 ;
    END
  END wd_in[525]
  PIN wd_in[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1081.325 0.070 1081.395 ;
    END
  END wd_in[526]
  PIN wd_in[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1081.465 0.070 1081.535 ;
    END
  END wd_in[527]
  PIN wd_in[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1081.605 0.070 1081.675 ;
    END
  END wd_in[528]
  PIN wd_in[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1081.745 0.070 1081.815 ;
    END
  END wd_in[529]
  PIN wd_in[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1081.885 0.070 1081.955 ;
    END
  END wd_in[530]
  PIN wd_in[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1082.025 0.070 1082.095 ;
    END
  END wd_in[531]
  PIN wd_in[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1082.165 0.070 1082.235 ;
    END
  END wd_in[532]
  PIN wd_in[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1082.305 0.070 1082.375 ;
    END
  END wd_in[533]
  PIN wd_in[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1082.445 0.070 1082.515 ;
    END
  END wd_in[534]
  PIN wd_in[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1082.585 0.070 1082.655 ;
    END
  END wd_in[535]
  PIN wd_in[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1082.725 0.070 1082.795 ;
    END
  END wd_in[536]
  PIN wd_in[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1082.865 0.070 1082.935 ;
    END
  END wd_in[537]
  PIN wd_in[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.005 0.070 1083.075 ;
    END
  END wd_in[538]
  PIN wd_in[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.145 0.070 1083.215 ;
    END
  END wd_in[539]
  PIN wd_in[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.285 0.070 1083.355 ;
    END
  END wd_in[540]
  PIN wd_in[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.425 0.070 1083.495 ;
    END
  END wd_in[541]
  PIN wd_in[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.565 0.070 1083.635 ;
    END
  END wd_in[542]
  PIN wd_in[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.705 0.070 1083.775 ;
    END
  END wd_in[543]
  PIN wd_in[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.845 0.070 1083.915 ;
    END
  END wd_in[544]
  PIN wd_in[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1083.985 0.070 1084.055 ;
    END
  END wd_in[545]
  PIN wd_in[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1084.125 0.070 1084.195 ;
    END
  END wd_in[546]
  PIN wd_in[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1084.265 0.070 1084.335 ;
    END
  END wd_in[547]
  PIN wd_in[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1084.405 0.070 1084.475 ;
    END
  END wd_in[548]
  PIN wd_in[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1084.545 0.070 1084.615 ;
    END
  END wd_in[549]
  PIN wd_in[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1084.685 0.070 1084.755 ;
    END
  END wd_in[550]
  PIN wd_in[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1084.825 0.070 1084.895 ;
    END
  END wd_in[551]
  PIN wd_in[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1084.965 0.070 1085.035 ;
    END
  END wd_in[552]
  PIN wd_in[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.105 0.070 1085.175 ;
    END
  END wd_in[553]
  PIN wd_in[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.245 0.070 1085.315 ;
    END
  END wd_in[554]
  PIN wd_in[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.385 0.070 1085.455 ;
    END
  END wd_in[555]
  PIN wd_in[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.525 0.070 1085.595 ;
    END
  END wd_in[556]
  PIN wd_in[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.665 0.070 1085.735 ;
    END
  END wd_in[557]
  PIN wd_in[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.805 0.070 1085.875 ;
    END
  END wd_in[558]
  PIN wd_in[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1085.945 0.070 1086.015 ;
    END
  END wd_in[559]
  PIN wd_in[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1086.085 0.070 1086.155 ;
    END
  END wd_in[560]
  PIN wd_in[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1086.225 0.070 1086.295 ;
    END
  END wd_in[561]
  PIN wd_in[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1086.365 0.070 1086.435 ;
    END
  END wd_in[562]
  PIN wd_in[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1086.505 0.070 1086.575 ;
    END
  END wd_in[563]
  PIN wd_in[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1086.645 0.070 1086.715 ;
    END
  END wd_in[564]
  PIN wd_in[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1086.785 0.070 1086.855 ;
    END
  END wd_in[565]
  PIN wd_in[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1086.925 0.070 1086.995 ;
    END
  END wd_in[566]
  PIN wd_in[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.065 0.070 1087.135 ;
    END
  END wd_in[567]
  PIN wd_in[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.205 0.070 1087.275 ;
    END
  END wd_in[568]
  PIN wd_in[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.345 0.070 1087.415 ;
    END
  END wd_in[569]
  PIN wd_in[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.485 0.070 1087.555 ;
    END
  END wd_in[570]
  PIN wd_in[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.625 0.070 1087.695 ;
    END
  END wd_in[571]
  PIN wd_in[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.765 0.070 1087.835 ;
    END
  END wd_in[572]
  PIN wd_in[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1087.905 0.070 1087.975 ;
    END
  END wd_in[573]
  PIN wd_in[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1088.045 0.070 1088.115 ;
    END
  END wd_in[574]
  PIN wd_in[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1088.185 0.070 1088.255 ;
    END
  END wd_in[575]
  PIN wd_in[576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1088.325 0.070 1088.395 ;
    END
  END wd_in[576]
  PIN wd_in[577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1088.465 0.070 1088.535 ;
    END
  END wd_in[577]
  PIN wd_in[578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1088.605 0.070 1088.675 ;
    END
  END wd_in[578]
  PIN wd_in[579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1088.745 0.070 1088.815 ;
    END
  END wd_in[579]
  PIN wd_in[580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1088.885 0.070 1088.955 ;
    END
  END wd_in[580]
  PIN wd_in[581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.025 0.070 1089.095 ;
    END
  END wd_in[581]
  PIN wd_in[582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.165 0.070 1089.235 ;
    END
  END wd_in[582]
  PIN wd_in[583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.305 0.070 1089.375 ;
    END
  END wd_in[583]
  PIN wd_in[584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.445 0.070 1089.515 ;
    END
  END wd_in[584]
  PIN wd_in[585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.585 0.070 1089.655 ;
    END
  END wd_in[585]
  PIN wd_in[586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.725 0.070 1089.795 ;
    END
  END wd_in[586]
  PIN wd_in[587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1089.865 0.070 1089.935 ;
    END
  END wd_in[587]
  PIN wd_in[588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.005 0.070 1090.075 ;
    END
  END wd_in[588]
  PIN wd_in[589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.145 0.070 1090.215 ;
    END
  END wd_in[589]
  PIN wd_in[590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.285 0.070 1090.355 ;
    END
  END wd_in[590]
  PIN wd_in[591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.425 0.070 1090.495 ;
    END
  END wd_in[591]
  PIN wd_in[592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.565 0.070 1090.635 ;
    END
  END wd_in[592]
  PIN wd_in[593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.705 0.070 1090.775 ;
    END
  END wd_in[593]
  PIN wd_in[594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.845 0.070 1090.915 ;
    END
  END wd_in[594]
  PIN wd_in[595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1090.985 0.070 1091.055 ;
    END
  END wd_in[595]
  PIN wd_in[596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1091.125 0.070 1091.195 ;
    END
  END wd_in[596]
  PIN wd_in[597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1091.265 0.070 1091.335 ;
    END
  END wd_in[597]
  PIN wd_in[598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1091.405 0.070 1091.475 ;
    END
  END wd_in[598]
  PIN wd_in[599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1091.545 0.070 1091.615 ;
    END
  END wd_in[599]
  PIN wd_in[600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1091.685 0.070 1091.755 ;
    END
  END wd_in[600]
  PIN wd_in[601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1091.825 0.070 1091.895 ;
    END
  END wd_in[601]
  PIN wd_in[602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1091.965 0.070 1092.035 ;
    END
  END wd_in[602]
  PIN wd_in[603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.105 0.070 1092.175 ;
    END
  END wd_in[603]
  PIN wd_in[604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.245 0.070 1092.315 ;
    END
  END wd_in[604]
  PIN wd_in[605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.385 0.070 1092.455 ;
    END
  END wd_in[605]
  PIN wd_in[606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.525 0.070 1092.595 ;
    END
  END wd_in[606]
  PIN wd_in[607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.665 0.070 1092.735 ;
    END
  END wd_in[607]
  PIN wd_in[608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.805 0.070 1092.875 ;
    END
  END wd_in[608]
  PIN wd_in[609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1092.945 0.070 1093.015 ;
    END
  END wd_in[609]
  PIN wd_in[610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1093.085 0.070 1093.155 ;
    END
  END wd_in[610]
  PIN wd_in[611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1093.225 0.070 1093.295 ;
    END
  END wd_in[611]
  PIN wd_in[612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1093.365 0.070 1093.435 ;
    END
  END wd_in[612]
  PIN wd_in[613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1093.505 0.070 1093.575 ;
    END
  END wd_in[613]
  PIN wd_in[614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1093.645 0.070 1093.715 ;
    END
  END wd_in[614]
  PIN wd_in[615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1093.785 0.070 1093.855 ;
    END
  END wd_in[615]
  PIN wd_in[616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1093.925 0.070 1093.995 ;
    END
  END wd_in[616]
  PIN wd_in[617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.065 0.070 1094.135 ;
    END
  END wd_in[617]
  PIN wd_in[618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.205 0.070 1094.275 ;
    END
  END wd_in[618]
  PIN wd_in[619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.345 0.070 1094.415 ;
    END
  END wd_in[619]
  PIN wd_in[620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.485 0.070 1094.555 ;
    END
  END wd_in[620]
  PIN wd_in[621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.625 0.070 1094.695 ;
    END
  END wd_in[621]
  PIN wd_in[622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.765 0.070 1094.835 ;
    END
  END wd_in[622]
  PIN wd_in[623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1094.905 0.070 1094.975 ;
    END
  END wd_in[623]
  PIN wd_in[624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1095.045 0.070 1095.115 ;
    END
  END wd_in[624]
  PIN wd_in[625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1095.185 0.070 1095.255 ;
    END
  END wd_in[625]
  PIN wd_in[626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1095.325 0.070 1095.395 ;
    END
  END wd_in[626]
  PIN wd_in[627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1095.465 0.070 1095.535 ;
    END
  END wd_in[627]
  PIN wd_in[628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1095.605 0.070 1095.675 ;
    END
  END wd_in[628]
  PIN wd_in[629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1095.745 0.070 1095.815 ;
    END
  END wd_in[629]
  PIN wd_in[630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1095.885 0.070 1095.955 ;
    END
  END wd_in[630]
  PIN wd_in[631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1096.025 0.070 1096.095 ;
    END
  END wd_in[631]
  PIN wd_in[632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1096.165 0.070 1096.235 ;
    END
  END wd_in[632]
  PIN wd_in[633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1096.305 0.070 1096.375 ;
    END
  END wd_in[633]
  PIN wd_in[634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1096.445 0.070 1096.515 ;
    END
  END wd_in[634]
  PIN wd_in[635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1096.585 0.070 1096.655 ;
    END
  END wd_in[635]
  PIN wd_in[636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1096.725 0.070 1096.795 ;
    END
  END wd_in[636]
  PIN wd_in[637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1096.865 0.070 1096.935 ;
    END
  END wd_in[637]
  PIN wd_in[638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.005 0.070 1097.075 ;
    END
  END wd_in[638]
  PIN wd_in[639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.145 0.070 1097.215 ;
    END
  END wd_in[639]
  PIN wd_in[640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.285 0.070 1097.355 ;
    END
  END wd_in[640]
  PIN wd_in[641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.425 0.070 1097.495 ;
    END
  END wd_in[641]
  PIN wd_in[642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.565 0.070 1097.635 ;
    END
  END wd_in[642]
  PIN wd_in[643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.705 0.070 1097.775 ;
    END
  END wd_in[643]
  PIN wd_in[644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.845 0.070 1097.915 ;
    END
  END wd_in[644]
  PIN wd_in[645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1097.985 0.070 1098.055 ;
    END
  END wd_in[645]
  PIN wd_in[646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1098.125 0.070 1098.195 ;
    END
  END wd_in[646]
  PIN wd_in[647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1098.265 0.070 1098.335 ;
    END
  END wd_in[647]
  PIN wd_in[648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1098.405 0.070 1098.475 ;
    END
  END wd_in[648]
  PIN wd_in[649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1098.545 0.070 1098.615 ;
    END
  END wd_in[649]
  PIN wd_in[650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1098.685 0.070 1098.755 ;
    END
  END wd_in[650]
  PIN wd_in[651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1098.825 0.070 1098.895 ;
    END
  END wd_in[651]
  PIN wd_in[652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1098.965 0.070 1099.035 ;
    END
  END wd_in[652]
  PIN wd_in[653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.105 0.070 1099.175 ;
    END
  END wd_in[653]
  PIN wd_in[654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.245 0.070 1099.315 ;
    END
  END wd_in[654]
  PIN wd_in[655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.385 0.070 1099.455 ;
    END
  END wd_in[655]
  PIN wd_in[656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.525 0.070 1099.595 ;
    END
  END wd_in[656]
  PIN wd_in[657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.665 0.070 1099.735 ;
    END
  END wd_in[657]
  PIN wd_in[658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.805 0.070 1099.875 ;
    END
  END wd_in[658]
  PIN wd_in[659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1099.945 0.070 1100.015 ;
    END
  END wd_in[659]
  PIN wd_in[660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.085 0.070 1100.155 ;
    END
  END wd_in[660]
  PIN wd_in[661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.225 0.070 1100.295 ;
    END
  END wd_in[661]
  PIN wd_in[662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.365 0.070 1100.435 ;
    END
  END wd_in[662]
  PIN wd_in[663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.505 0.070 1100.575 ;
    END
  END wd_in[663]
  PIN wd_in[664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.645 0.070 1100.715 ;
    END
  END wd_in[664]
  PIN wd_in[665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.785 0.070 1100.855 ;
    END
  END wd_in[665]
  PIN wd_in[666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1100.925 0.070 1100.995 ;
    END
  END wd_in[666]
  PIN wd_in[667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.065 0.070 1101.135 ;
    END
  END wd_in[667]
  PIN wd_in[668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.205 0.070 1101.275 ;
    END
  END wd_in[668]
  PIN wd_in[669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.345 0.070 1101.415 ;
    END
  END wd_in[669]
  PIN wd_in[670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.485 0.070 1101.555 ;
    END
  END wd_in[670]
  PIN wd_in[671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.625 0.070 1101.695 ;
    END
  END wd_in[671]
  PIN wd_in[672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.765 0.070 1101.835 ;
    END
  END wd_in[672]
  PIN wd_in[673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1101.905 0.070 1101.975 ;
    END
  END wd_in[673]
  PIN wd_in[674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1102.045 0.070 1102.115 ;
    END
  END wd_in[674]
  PIN wd_in[675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1102.185 0.070 1102.255 ;
    END
  END wd_in[675]
  PIN wd_in[676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1102.325 0.070 1102.395 ;
    END
  END wd_in[676]
  PIN wd_in[677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1102.465 0.070 1102.535 ;
    END
  END wd_in[677]
  PIN wd_in[678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1102.605 0.070 1102.675 ;
    END
  END wd_in[678]
  PIN wd_in[679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1102.745 0.070 1102.815 ;
    END
  END wd_in[679]
  PIN wd_in[680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1102.885 0.070 1102.955 ;
    END
  END wd_in[680]
  PIN wd_in[681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1103.025 0.070 1103.095 ;
    END
  END wd_in[681]
  PIN wd_in[682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1103.165 0.070 1103.235 ;
    END
  END wd_in[682]
  PIN wd_in[683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1103.305 0.070 1103.375 ;
    END
  END wd_in[683]
  PIN wd_in[684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1103.445 0.070 1103.515 ;
    END
  END wd_in[684]
  PIN wd_in[685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1103.585 0.070 1103.655 ;
    END
  END wd_in[685]
  PIN wd_in[686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1103.725 0.070 1103.795 ;
    END
  END wd_in[686]
  PIN wd_in[687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1103.865 0.070 1103.935 ;
    END
  END wd_in[687]
  PIN wd_in[688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.005 0.070 1104.075 ;
    END
  END wd_in[688]
  PIN wd_in[689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.145 0.070 1104.215 ;
    END
  END wd_in[689]
  PIN wd_in[690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.285 0.070 1104.355 ;
    END
  END wd_in[690]
  PIN wd_in[691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.425 0.070 1104.495 ;
    END
  END wd_in[691]
  PIN wd_in[692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.565 0.070 1104.635 ;
    END
  END wd_in[692]
  PIN wd_in[693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.705 0.070 1104.775 ;
    END
  END wd_in[693]
  PIN wd_in[694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.845 0.070 1104.915 ;
    END
  END wd_in[694]
  PIN wd_in[695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1104.985 0.070 1105.055 ;
    END
  END wd_in[695]
  PIN wd_in[696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1105.125 0.070 1105.195 ;
    END
  END wd_in[696]
  PIN wd_in[697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1105.265 0.070 1105.335 ;
    END
  END wd_in[697]
  PIN wd_in[698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1105.405 0.070 1105.475 ;
    END
  END wd_in[698]
  PIN wd_in[699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1105.545 0.070 1105.615 ;
    END
  END wd_in[699]
  PIN wd_in[700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1105.685 0.070 1105.755 ;
    END
  END wd_in[700]
  PIN wd_in[701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1105.825 0.070 1105.895 ;
    END
  END wd_in[701]
  PIN wd_in[702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1105.965 0.070 1106.035 ;
    END
  END wd_in[702]
  PIN wd_in[703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.105 0.070 1106.175 ;
    END
  END wd_in[703]
  PIN wd_in[704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.245 0.070 1106.315 ;
    END
  END wd_in[704]
  PIN wd_in[705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.385 0.070 1106.455 ;
    END
  END wd_in[705]
  PIN wd_in[706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.525 0.070 1106.595 ;
    END
  END wd_in[706]
  PIN wd_in[707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.665 0.070 1106.735 ;
    END
  END wd_in[707]
  PIN wd_in[708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.805 0.070 1106.875 ;
    END
  END wd_in[708]
  PIN wd_in[709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1106.945 0.070 1107.015 ;
    END
  END wd_in[709]
  PIN wd_in[710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1107.085 0.070 1107.155 ;
    END
  END wd_in[710]
  PIN wd_in[711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1107.225 0.070 1107.295 ;
    END
  END wd_in[711]
  PIN wd_in[712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1107.365 0.070 1107.435 ;
    END
  END wd_in[712]
  PIN wd_in[713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1107.505 0.070 1107.575 ;
    END
  END wd_in[713]
  PIN wd_in[714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1107.645 0.070 1107.715 ;
    END
  END wd_in[714]
  PIN wd_in[715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1107.785 0.070 1107.855 ;
    END
  END wd_in[715]
  PIN wd_in[716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1107.925 0.070 1107.995 ;
    END
  END wd_in[716]
  PIN wd_in[717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.065 0.070 1108.135 ;
    END
  END wd_in[717]
  PIN wd_in[718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.205 0.070 1108.275 ;
    END
  END wd_in[718]
  PIN wd_in[719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.345 0.070 1108.415 ;
    END
  END wd_in[719]
  PIN wd_in[720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.485 0.070 1108.555 ;
    END
  END wd_in[720]
  PIN wd_in[721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.625 0.070 1108.695 ;
    END
  END wd_in[721]
  PIN wd_in[722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.765 0.070 1108.835 ;
    END
  END wd_in[722]
  PIN wd_in[723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1108.905 0.070 1108.975 ;
    END
  END wd_in[723]
  PIN wd_in[724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1109.045 0.070 1109.115 ;
    END
  END wd_in[724]
  PIN wd_in[725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1109.185 0.070 1109.255 ;
    END
  END wd_in[725]
  PIN wd_in[726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1109.325 0.070 1109.395 ;
    END
  END wd_in[726]
  PIN wd_in[727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1109.465 0.070 1109.535 ;
    END
  END wd_in[727]
  PIN wd_in[728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1109.605 0.070 1109.675 ;
    END
  END wd_in[728]
  PIN wd_in[729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1109.745 0.070 1109.815 ;
    END
  END wd_in[729]
  PIN wd_in[730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1109.885 0.070 1109.955 ;
    END
  END wd_in[730]
  PIN wd_in[731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1110.025 0.070 1110.095 ;
    END
  END wd_in[731]
  PIN wd_in[732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1110.165 0.070 1110.235 ;
    END
  END wd_in[732]
  PIN wd_in[733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1110.305 0.070 1110.375 ;
    END
  END wd_in[733]
  PIN wd_in[734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1110.445 0.070 1110.515 ;
    END
  END wd_in[734]
  PIN wd_in[735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1110.585 0.070 1110.655 ;
    END
  END wd_in[735]
  PIN wd_in[736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1110.725 0.070 1110.795 ;
    END
  END wd_in[736]
  PIN wd_in[737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1110.865 0.070 1110.935 ;
    END
  END wd_in[737]
  PIN wd_in[738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.005 0.070 1111.075 ;
    END
  END wd_in[738]
  PIN wd_in[739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.145 0.070 1111.215 ;
    END
  END wd_in[739]
  PIN wd_in[740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.285 0.070 1111.355 ;
    END
  END wd_in[740]
  PIN wd_in[741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.425 0.070 1111.495 ;
    END
  END wd_in[741]
  PIN wd_in[742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.565 0.070 1111.635 ;
    END
  END wd_in[742]
  PIN wd_in[743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.705 0.070 1111.775 ;
    END
  END wd_in[743]
  PIN wd_in[744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.845 0.070 1111.915 ;
    END
  END wd_in[744]
  PIN wd_in[745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1111.985 0.070 1112.055 ;
    END
  END wd_in[745]
  PIN wd_in[746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1112.125 0.070 1112.195 ;
    END
  END wd_in[746]
  PIN wd_in[747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1112.265 0.070 1112.335 ;
    END
  END wd_in[747]
  PIN wd_in[748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1112.405 0.070 1112.475 ;
    END
  END wd_in[748]
  PIN wd_in[749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1112.545 0.070 1112.615 ;
    END
  END wd_in[749]
  PIN wd_in[750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1112.685 0.070 1112.755 ;
    END
  END wd_in[750]
  PIN wd_in[751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1112.825 0.070 1112.895 ;
    END
  END wd_in[751]
  PIN wd_in[752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1112.965 0.070 1113.035 ;
    END
  END wd_in[752]
  PIN wd_in[753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.105 0.070 1113.175 ;
    END
  END wd_in[753]
  PIN wd_in[754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.245 0.070 1113.315 ;
    END
  END wd_in[754]
  PIN wd_in[755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.385 0.070 1113.455 ;
    END
  END wd_in[755]
  PIN wd_in[756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.525 0.070 1113.595 ;
    END
  END wd_in[756]
  PIN wd_in[757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.665 0.070 1113.735 ;
    END
  END wd_in[757]
  PIN wd_in[758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.805 0.070 1113.875 ;
    END
  END wd_in[758]
  PIN wd_in[759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1113.945 0.070 1114.015 ;
    END
  END wd_in[759]
  PIN wd_in[760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1114.085 0.070 1114.155 ;
    END
  END wd_in[760]
  PIN wd_in[761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1114.225 0.070 1114.295 ;
    END
  END wd_in[761]
  PIN wd_in[762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1114.365 0.070 1114.435 ;
    END
  END wd_in[762]
  PIN wd_in[763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1114.505 0.070 1114.575 ;
    END
  END wd_in[763]
  PIN wd_in[764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1114.645 0.070 1114.715 ;
    END
  END wd_in[764]
  PIN wd_in[765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1114.785 0.070 1114.855 ;
    END
  END wd_in[765]
  PIN wd_in[766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1114.925 0.070 1114.995 ;
    END
  END wd_in[766]
  PIN wd_in[767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.065 0.070 1115.135 ;
    END
  END wd_in[767]
  PIN wd_in[768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.205 0.070 1115.275 ;
    END
  END wd_in[768]
  PIN wd_in[769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.345 0.070 1115.415 ;
    END
  END wd_in[769]
  PIN wd_in[770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.485 0.070 1115.555 ;
    END
  END wd_in[770]
  PIN wd_in[771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.625 0.070 1115.695 ;
    END
  END wd_in[771]
  PIN wd_in[772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.765 0.070 1115.835 ;
    END
  END wd_in[772]
  PIN wd_in[773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1115.905 0.070 1115.975 ;
    END
  END wd_in[773]
  PIN wd_in[774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1116.045 0.070 1116.115 ;
    END
  END wd_in[774]
  PIN wd_in[775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1116.185 0.070 1116.255 ;
    END
  END wd_in[775]
  PIN wd_in[776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1116.325 0.070 1116.395 ;
    END
  END wd_in[776]
  PIN wd_in[777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1116.465 0.070 1116.535 ;
    END
  END wd_in[777]
  PIN wd_in[778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1116.605 0.070 1116.675 ;
    END
  END wd_in[778]
  PIN wd_in[779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1116.745 0.070 1116.815 ;
    END
  END wd_in[779]
  PIN wd_in[780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1116.885 0.070 1116.955 ;
    END
  END wd_in[780]
  PIN wd_in[781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1117.025 0.070 1117.095 ;
    END
  END wd_in[781]
  PIN wd_in[782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1117.165 0.070 1117.235 ;
    END
  END wd_in[782]
  PIN wd_in[783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1117.305 0.070 1117.375 ;
    END
  END wd_in[783]
  PIN wd_in[784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1117.445 0.070 1117.515 ;
    END
  END wd_in[784]
  PIN wd_in[785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1117.585 0.070 1117.655 ;
    END
  END wd_in[785]
  PIN wd_in[786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1117.725 0.070 1117.795 ;
    END
  END wd_in[786]
  PIN wd_in[787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1117.865 0.070 1117.935 ;
    END
  END wd_in[787]
  PIN wd_in[788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.005 0.070 1118.075 ;
    END
  END wd_in[788]
  PIN wd_in[789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.145 0.070 1118.215 ;
    END
  END wd_in[789]
  PIN wd_in[790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.285 0.070 1118.355 ;
    END
  END wd_in[790]
  PIN wd_in[791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.425 0.070 1118.495 ;
    END
  END wd_in[791]
  PIN wd_in[792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.565 0.070 1118.635 ;
    END
  END wd_in[792]
  PIN wd_in[793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.705 0.070 1118.775 ;
    END
  END wd_in[793]
  PIN wd_in[794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.845 0.070 1118.915 ;
    END
  END wd_in[794]
  PIN wd_in[795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1118.985 0.070 1119.055 ;
    END
  END wd_in[795]
  PIN wd_in[796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1119.125 0.070 1119.195 ;
    END
  END wd_in[796]
  PIN wd_in[797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1119.265 0.070 1119.335 ;
    END
  END wd_in[797]
  PIN wd_in[798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1119.405 0.070 1119.475 ;
    END
  END wd_in[798]
  PIN wd_in[799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1119.545 0.070 1119.615 ;
    END
  END wd_in[799]
  PIN wd_in[800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1119.685 0.070 1119.755 ;
    END
  END wd_in[800]
  PIN wd_in[801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1119.825 0.070 1119.895 ;
    END
  END wd_in[801]
  PIN wd_in[802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1119.965 0.070 1120.035 ;
    END
  END wd_in[802]
  PIN wd_in[803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.105 0.070 1120.175 ;
    END
  END wd_in[803]
  PIN wd_in[804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.245 0.070 1120.315 ;
    END
  END wd_in[804]
  PIN wd_in[805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.385 0.070 1120.455 ;
    END
  END wd_in[805]
  PIN wd_in[806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.525 0.070 1120.595 ;
    END
  END wd_in[806]
  PIN wd_in[807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.665 0.070 1120.735 ;
    END
  END wd_in[807]
  PIN wd_in[808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.805 0.070 1120.875 ;
    END
  END wd_in[808]
  PIN wd_in[809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1120.945 0.070 1121.015 ;
    END
  END wd_in[809]
  PIN wd_in[810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.085 0.070 1121.155 ;
    END
  END wd_in[810]
  PIN wd_in[811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.225 0.070 1121.295 ;
    END
  END wd_in[811]
  PIN wd_in[812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.365 0.070 1121.435 ;
    END
  END wd_in[812]
  PIN wd_in[813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.505 0.070 1121.575 ;
    END
  END wd_in[813]
  PIN wd_in[814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.645 0.070 1121.715 ;
    END
  END wd_in[814]
  PIN wd_in[815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.785 0.070 1121.855 ;
    END
  END wd_in[815]
  PIN wd_in[816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1121.925 0.070 1121.995 ;
    END
  END wd_in[816]
  PIN wd_in[817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.065 0.070 1122.135 ;
    END
  END wd_in[817]
  PIN wd_in[818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.205 0.070 1122.275 ;
    END
  END wd_in[818]
  PIN wd_in[819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.345 0.070 1122.415 ;
    END
  END wd_in[819]
  PIN wd_in[820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.485 0.070 1122.555 ;
    END
  END wd_in[820]
  PIN wd_in[821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.625 0.070 1122.695 ;
    END
  END wd_in[821]
  PIN wd_in[822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.765 0.070 1122.835 ;
    END
  END wd_in[822]
  PIN wd_in[823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1122.905 0.070 1122.975 ;
    END
  END wd_in[823]
  PIN wd_in[824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1123.045 0.070 1123.115 ;
    END
  END wd_in[824]
  PIN wd_in[825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1123.185 0.070 1123.255 ;
    END
  END wd_in[825]
  PIN wd_in[826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1123.325 0.070 1123.395 ;
    END
  END wd_in[826]
  PIN wd_in[827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1123.465 0.070 1123.535 ;
    END
  END wd_in[827]
  PIN wd_in[828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1123.605 0.070 1123.675 ;
    END
  END wd_in[828]
  PIN wd_in[829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1123.745 0.070 1123.815 ;
    END
  END wd_in[829]
  PIN wd_in[830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1123.885 0.070 1123.955 ;
    END
  END wd_in[830]
  PIN wd_in[831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1124.025 0.070 1124.095 ;
    END
  END wd_in[831]
  PIN wd_in[832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1124.165 0.070 1124.235 ;
    END
  END wd_in[832]
  PIN wd_in[833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1124.305 0.070 1124.375 ;
    END
  END wd_in[833]
  PIN wd_in[834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1124.445 0.070 1124.515 ;
    END
  END wd_in[834]
  PIN wd_in[835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1124.585 0.070 1124.655 ;
    END
  END wd_in[835]
  PIN wd_in[836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1124.725 0.070 1124.795 ;
    END
  END wd_in[836]
  PIN wd_in[837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1124.865 0.070 1124.935 ;
    END
  END wd_in[837]
  PIN wd_in[838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.005 0.070 1125.075 ;
    END
  END wd_in[838]
  PIN wd_in[839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.145 0.070 1125.215 ;
    END
  END wd_in[839]
  PIN wd_in[840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.285 0.070 1125.355 ;
    END
  END wd_in[840]
  PIN wd_in[841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.425 0.070 1125.495 ;
    END
  END wd_in[841]
  PIN wd_in[842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.565 0.070 1125.635 ;
    END
  END wd_in[842]
  PIN wd_in[843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.705 0.070 1125.775 ;
    END
  END wd_in[843]
  PIN wd_in[844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.845 0.070 1125.915 ;
    END
  END wd_in[844]
  PIN wd_in[845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1125.985 0.070 1126.055 ;
    END
  END wd_in[845]
  PIN wd_in[846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1126.125 0.070 1126.195 ;
    END
  END wd_in[846]
  PIN wd_in[847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1126.265 0.070 1126.335 ;
    END
  END wd_in[847]
  PIN wd_in[848]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1126.405 0.070 1126.475 ;
    END
  END wd_in[848]
  PIN wd_in[849]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1126.545 0.070 1126.615 ;
    END
  END wd_in[849]
  PIN wd_in[850]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1126.685 0.070 1126.755 ;
    END
  END wd_in[850]
  PIN wd_in[851]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1126.825 0.070 1126.895 ;
    END
  END wd_in[851]
  PIN wd_in[852]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1126.965 0.070 1127.035 ;
    END
  END wd_in[852]
  PIN wd_in[853]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.105 0.070 1127.175 ;
    END
  END wd_in[853]
  PIN wd_in[854]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.245 0.070 1127.315 ;
    END
  END wd_in[854]
  PIN wd_in[855]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.385 0.070 1127.455 ;
    END
  END wd_in[855]
  PIN wd_in[856]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.525 0.070 1127.595 ;
    END
  END wd_in[856]
  PIN wd_in[857]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.665 0.070 1127.735 ;
    END
  END wd_in[857]
  PIN wd_in[858]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.805 0.070 1127.875 ;
    END
  END wd_in[858]
  PIN wd_in[859]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1127.945 0.070 1128.015 ;
    END
  END wd_in[859]
  PIN wd_in[860]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1128.085 0.070 1128.155 ;
    END
  END wd_in[860]
  PIN wd_in[861]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1128.225 0.070 1128.295 ;
    END
  END wd_in[861]
  PIN wd_in[862]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1128.365 0.070 1128.435 ;
    END
  END wd_in[862]
  PIN wd_in[863]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1128.505 0.070 1128.575 ;
    END
  END wd_in[863]
  PIN wd_in[864]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1128.645 0.070 1128.715 ;
    END
  END wd_in[864]
  PIN wd_in[865]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1128.785 0.070 1128.855 ;
    END
  END wd_in[865]
  PIN wd_in[866]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1128.925 0.070 1128.995 ;
    END
  END wd_in[866]
  PIN wd_in[867]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.065 0.070 1129.135 ;
    END
  END wd_in[867]
  PIN wd_in[868]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.205 0.070 1129.275 ;
    END
  END wd_in[868]
  PIN wd_in[869]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.345 0.070 1129.415 ;
    END
  END wd_in[869]
  PIN wd_in[870]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.485 0.070 1129.555 ;
    END
  END wd_in[870]
  PIN wd_in[871]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.625 0.070 1129.695 ;
    END
  END wd_in[871]
  PIN wd_in[872]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.765 0.070 1129.835 ;
    END
  END wd_in[872]
  PIN wd_in[873]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1129.905 0.070 1129.975 ;
    END
  END wd_in[873]
  PIN wd_in[874]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1130.045 0.070 1130.115 ;
    END
  END wd_in[874]
  PIN wd_in[875]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1130.185 0.070 1130.255 ;
    END
  END wd_in[875]
  PIN wd_in[876]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1130.325 0.070 1130.395 ;
    END
  END wd_in[876]
  PIN wd_in[877]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1130.465 0.070 1130.535 ;
    END
  END wd_in[877]
  PIN wd_in[878]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1130.605 0.070 1130.675 ;
    END
  END wd_in[878]
  PIN wd_in[879]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1130.745 0.070 1130.815 ;
    END
  END wd_in[879]
  PIN wd_in[880]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1130.885 0.070 1130.955 ;
    END
  END wd_in[880]
  PIN wd_in[881]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1131.025 0.070 1131.095 ;
    END
  END wd_in[881]
  PIN wd_in[882]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1131.165 0.070 1131.235 ;
    END
  END wd_in[882]
  PIN wd_in[883]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1131.305 0.070 1131.375 ;
    END
  END wd_in[883]
  PIN wd_in[884]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1131.445 0.070 1131.515 ;
    END
  END wd_in[884]
  PIN wd_in[885]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1131.585 0.070 1131.655 ;
    END
  END wd_in[885]
  PIN wd_in[886]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1131.725 0.070 1131.795 ;
    END
  END wd_in[886]
  PIN wd_in[887]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1131.865 0.070 1131.935 ;
    END
  END wd_in[887]
  PIN wd_in[888]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.005 0.070 1132.075 ;
    END
  END wd_in[888]
  PIN wd_in[889]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.145 0.070 1132.215 ;
    END
  END wd_in[889]
  PIN wd_in[890]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.285 0.070 1132.355 ;
    END
  END wd_in[890]
  PIN wd_in[891]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.425 0.070 1132.495 ;
    END
  END wd_in[891]
  PIN wd_in[892]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.565 0.070 1132.635 ;
    END
  END wd_in[892]
  PIN wd_in[893]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.705 0.070 1132.775 ;
    END
  END wd_in[893]
  PIN wd_in[894]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.845 0.070 1132.915 ;
    END
  END wd_in[894]
  PIN wd_in[895]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1132.985 0.070 1133.055 ;
    END
  END wd_in[895]
  PIN wd_in[896]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1133.125 0.070 1133.195 ;
    END
  END wd_in[896]
  PIN wd_in[897]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1133.265 0.070 1133.335 ;
    END
  END wd_in[897]
  PIN wd_in[898]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1133.405 0.070 1133.475 ;
    END
  END wd_in[898]
  PIN wd_in[899]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1133.545 0.070 1133.615 ;
    END
  END wd_in[899]
  PIN wd_in[900]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1133.685 0.070 1133.755 ;
    END
  END wd_in[900]
  PIN wd_in[901]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1133.825 0.070 1133.895 ;
    END
  END wd_in[901]
  PIN wd_in[902]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1133.965 0.070 1134.035 ;
    END
  END wd_in[902]
  PIN wd_in[903]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.105 0.070 1134.175 ;
    END
  END wd_in[903]
  PIN wd_in[904]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.245 0.070 1134.315 ;
    END
  END wd_in[904]
  PIN wd_in[905]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.385 0.070 1134.455 ;
    END
  END wd_in[905]
  PIN wd_in[906]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.525 0.070 1134.595 ;
    END
  END wd_in[906]
  PIN wd_in[907]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.665 0.070 1134.735 ;
    END
  END wd_in[907]
  PIN wd_in[908]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.805 0.070 1134.875 ;
    END
  END wd_in[908]
  PIN wd_in[909]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1134.945 0.070 1135.015 ;
    END
  END wd_in[909]
  PIN wd_in[910]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1135.085 0.070 1135.155 ;
    END
  END wd_in[910]
  PIN wd_in[911]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1135.225 0.070 1135.295 ;
    END
  END wd_in[911]
  PIN wd_in[912]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1135.365 0.070 1135.435 ;
    END
  END wd_in[912]
  PIN wd_in[913]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1135.505 0.070 1135.575 ;
    END
  END wd_in[913]
  PIN wd_in[914]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1135.645 0.070 1135.715 ;
    END
  END wd_in[914]
  PIN wd_in[915]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1135.785 0.070 1135.855 ;
    END
  END wd_in[915]
  PIN wd_in[916]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1135.925 0.070 1135.995 ;
    END
  END wd_in[916]
  PIN wd_in[917]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.065 0.070 1136.135 ;
    END
  END wd_in[917]
  PIN wd_in[918]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.205 0.070 1136.275 ;
    END
  END wd_in[918]
  PIN wd_in[919]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.345 0.070 1136.415 ;
    END
  END wd_in[919]
  PIN wd_in[920]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.485 0.070 1136.555 ;
    END
  END wd_in[920]
  PIN wd_in[921]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.625 0.070 1136.695 ;
    END
  END wd_in[921]
  PIN wd_in[922]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.765 0.070 1136.835 ;
    END
  END wd_in[922]
  PIN wd_in[923]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1136.905 0.070 1136.975 ;
    END
  END wd_in[923]
  PIN wd_in[924]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1137.045 0.070 1137.115 ;
    END
  END wd_in[924]
  PIN wd_in[925]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1137.185 0.070 1137.255 ;
    END
  END wd_in[925]
  PIN wd_in[926]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1137.325 0.070 1137.395 ;
    END
  END wd_in[926]
  PIN wd_in[927]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1137.465 0.070 1137.535 ;
    END
  END wd_in[927]
  PIN wd_in[928]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1137.605 0.070 1137.675 ;
    END
  END wd_in[928]
  PIN wd_in[929]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1137.745 0.070 1137.815 ;
    END
  END wd_in[929]
  PIN wd_in[930]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1137.885 0.070 1137.955 ;
    END
  END wd_in[930]
  PIN wd_in[931]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1138.025 0.070 1138.095 ;
    END
  END wd_in[931]
  PIN wd_in[932]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1138.165 0.070 1138.235 ;
    END
  END wd_in[932]
  PIN wd_in[933]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1138.305 0.070 1138.375 ;
    END
  END wd_in[933]
  PIN wd_in[934]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1138.445 0.070 1138.515 ;
    END
  END wd_in[934]
  PIN wd_in[935]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1138.585 0.070 1138.655 ;
    END
  END wd_in[935]
  PIN wd_in[936]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1138.725 0.070 1138.795 ;
    END
  END wd_in[936]
  PIN wd_in[937]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1138.865 0.070 1138.935 ;
    END
  END wd_in[937]
  PIN wd_in[938]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.005 0.070 1139.075 ;
    END
  END wd_in[938]
  PIN wd_in[939]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.145 0.070 1139.215 ;
    END
  END wd_in[939]
  PIN wd_in[940]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.285 0.070 1139.355 ;
    END
  END wd_in[940]
  PIN wd_in[941]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.425 0.070 1139.495 ;
    END
  END wd_in[941]
  PIN wd_in[942]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.565 0.070 1139.635 ;
    END
  END wd_in[942]
  PIN wd_in[943]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.705 0.070 1139.775 ;
    END
  END wd_in[943]
  PIN wd_in[944]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.845 0.070 1139.915 ;
    END
  END wd_in[944]
  PIN wd_in[945]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1139.985 0.070 1140.055 ;
    END
  END wd_in[945]
  PIN wd_in[946]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1140.125 0.070 1140.195 ;
    END
  END wd_in[946]
  PIN wd_in[947]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1140.265 0.070 1140.335 ;
    END
  END wd_in[947]
  PIN wd_in[948]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1140.405 0.070 1140.475 ;
    END
  END wd_in[948]
  PIN wd_in[949]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1140.545 0.070 1140.615 ;
    END
  END wd_in[949]
  PIN wd_in[950]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1140.685 0.070 1140.755 ;
    END
  END wd_in[950]
  PIN wd_in[951]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1140.825 0.070 1140.895 ;
    END
  END wd_in[951]
  PIN wd_in[952]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1140.965 0.070 1141.035 ;
    END
  END wd_in[952]
  PIN wd_in[953]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.105 0.070 1141.175 ;
    END
  END wd_in[953]
  PIN wd_in[954]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.245 0.070 1141.315 ;
    END
  END wd_in[954]
  PIN wd_in[955]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.385 0.070 1141.455 ;
    END
  END wd_in[955]
  PIN wd_in[956]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.525 0.070 1141.595 ;
    END
  END wd_in[956]
  PIN wd_in[957]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.665 0.070 1141.735 ;
    END
  END wd_in[957]
  PIN wd_in[958]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.805 0.070 1141.875 ;
    END
  END wd_in[958]
  PIN wd_in[959]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1141.945 0.070 1142.015 ;
    END
  END wd_in[959]
  PIN wd_in[960]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1142.085 0.070 1142.155 ;
    END
  END wd_in[960]
  PIN wd_in[961]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1142.225 0.070 1142.295 ;
    END
  END wd_in[961]
  PIN wd_in[962]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1142.365 0.070 1142.435 ;
    END
  END wd_in[962]
  PIN wd_in[963]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1142.505 0.070 1142.575 ;
    END
  END wd_in[963]
  PIN wd_in[964]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1142.645 0.070 1142.715 ;
    END
  END wd_in[964]
  PIN wd_in[965]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1142.785 0.070 1142.855 ;
    END
  END wd_in[965]
  PIN wd_in[966]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1142.925 0.070 1142.995 ;
    END
  END wd_in[966]
  PIN wd_in[967]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.065 0.070 1143.135 ;
    END
  END wd_in[967]
  PIN wd_in[968]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.205 0.070 1143.275 ;
    END
  END wd_in[968]
  PIN wd_in[969]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.345 0.070 1143.415 ;
    END
  END wd_in[969]
  PIN wd_in[970]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.485 0.070 1143.555 ;
    END
  END wd_in[970]
  PIN wd_in[971]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.625 0.070 1143.695 ;
    END
  END wd_in[971]
  PIN wd_in[972]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.765 0.070 1143.835 ;
    END
  END wd_in[972]
  PIN wd_in[973]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1143.905 0.070 1143.975 ;
    END
  END wd_in[973]
  PIN wd_in[974]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1144.045 0.070 1144.115 ;
    END
  END wd_in[974]
  PIN wd_in[975]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1144.185 0.070 1144.255 ;
    END
  END wd_in[975]
  PIN wd_in[976]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1144.325 0.070 1144.395 ;
    END
  END wd_in[976]
  PIN wd_in[977]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1144.465 0.070 1144.535 ;
    END
  END wd_in[977]
  PIN wd_in[978]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1144.605 0.070 1144.675 ;
    END
  END wd_in[978]
  PIN wd_in[979]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1144.745 0.070 1144.815 ;
    END
  END wd_in[979]
  PIN wd_in[980]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1144.885 0.070 1144.955 ;
    END
  END wd_in[980]
  PIN wd_in[981]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1145.025 0.070 1145.095 ;
    END
  END wd_in[981]
  PIN wd_in[982]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1145.165 0.070 1145.235 ;
    END
  END wd_in[982]
  PIN wd_in[983]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1145.305 0.070 1145.375 ;
    END
  END wd_in[983]
  PIN wd_in[984]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1145.445 0.070 1145.515 ;
    END
  END wd_in[984]
  PIN wd_in[985]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1145.585 0.070 1145.655 ;
    END
  END wd_in[985]
  PIN wd_in[986]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1145.725 0.070 1145.795 ;
    END
  END wd_in[986]
  PIN wd_in[987]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1145.865 0.070 1145.935 ;
    END
  END wd_in[987]
  PIN wd_in[988]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.005 0.070 1146.075 ;
    END
  END wd_in[988]
  PIN wd_in[989]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.145 0.070 1146.215 ;
    END
  END wd_in[989]
  PIN wd_in[990]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.285 0.070 1146.355 ;
    END
  END wd_in[990]
  PIN wd_in[991]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.425 0.070 1146.495 ;
    END
  END wd_in[991]
  PIN wd_in[992]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.565 0.070 1146.635 ;
    END
  END wd_in[992]
  PIN wd_in[993]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.705 0.070 1146.775 ;
    END
  END wd_in[993]
  PIN wd_in[994]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.845 0.070 1146.915 ;
    END
  END wd_in[994]
  PIN wd_in[995]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1146.985 0.070 1147.055 ;
    END
  END wd_in[995]
  PIN wd_in[996]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1147.125 0.070 1147.195 ;
    END
  END wd_in[996]
  PIN wd_in[997]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1147.265 0.070 1147.335 ;
    END
  END wd_in[997]
  PIN wd_in[998]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1147.405 0.070 1147.475 ;
    END
  END wd_in[998]
  PIN wd_in[999]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1147.545 0.070 1147.615 ;
    END
  END wd_in[999]
  PIN wd_in[1000]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1147.685 0.070 1147.755 ;
    END
  END wd_in[1000]
  PIN wd_in[1001]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1147.825 0.070 1147.895 ;
    END
  END wd_in[1001]
  PIN wd_in[1002]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1147.965 0.070 1148.035 ;
    END
  END wd_in[1002]
  PIN wd_in[1003]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.105 0.070 1148.175 ;
    END
  END wd_in[1003]
  PIN wd_in[1004]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.245 0.070 1148.315 ;
    END
  END wd_in[1004]
  PIN wd_in[1005]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.385 0.070 1148.455 ;
    END
  END wd_in[1005]
  PIN wd_in[1006]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.525 0.070 1148.595 ;
    END
  END wd_in[1006]
  PIN wd_in[1007]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.665 0.070 1148.735 ;
    END
  END wd_in[1007]
  PIN wd_in[1008]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.805 0.070 1148.875 ;
    END
  END wd_in[1008]
  PIN wd_in[1009]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1148.945 0.070 1149.015 ;
    END
  END wd_in[1009]
  PIN wd_in[1010]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1149.085 0.070 1149.155 ;
    END
  END wd_in[1010]
  PIN wd_in[1011]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1149.225 0.070 1149.295 ;
    END
  END wd_in[1011]
  PIN wd_in[1012]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1149.365 0.070 1149.435 ;
    END
  END wd_in[1012]
  PIN wd_in[1013]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1149.505 0.070 1149.575 ;
    END
  END wd_in[1013]
  PIN wd_in[1014]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1149.645 0.070 1149.715 ;
    END
  END wd_in[1014]
  PIN wd_in[1015]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1149.785 0.070 1149.855 ;
    END
  END wd_in[1015]
  PIN wd_in[1016]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1149.925 0.070 1149.995 ;
    END
  END wd_in[1016]
  PIN wd_in[1017]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.065 0.070 1150.135 ;
    END
  END wd_in[1017]
  PIN wd_in[1018]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.205 0.070 1150.275 ;
    END
  END wd_in[1018]
  PIN wd_in[1019]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.345 0.070 1150.415 ;
    END
  END wd_in[1019]
  PIN wd_in[1020]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.485 0.070 1150.555 ;
    END
  END wd_in[1020]
  PIN wd_in[1021]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.625 0.070 1150.695 ;
    END
  END wd_in[1021]
  PIN wd_in[1022]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.765 0.070 1150.835 ;
    END
  END wd_in[1022]
  PIN wd_in[1023]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1150.905 0.070 1150.975 ;
    END
  END wd_in[1023]
  PIN wd_in[1024]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1151.045 0.070 1151.115 ;
    END
  END wd_in[1024]
  PIN wd_in[1025]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1151.185 0.070 1151.255 ;
    END
  END wd_in[1025]
  PIN wd_in[1026]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1151.325 0.070 1151.395 ;
    END
  END wd_in[1026]
  PIN wd_in[1027]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1151.465 0.070 1151.535 ;
    END
  END wd_in[1027]
  PIN wd_in[1028]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1151.605 0.070 1151.675 ;
    END
  END wd_in[1028]
  PIN wd_in[1029]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1151.745 0.070 1151.815 ;
    END
  END wd_in[1029]
  PIN wd_in[1030]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1151.885 0.070 1151.955 ;
    END
  END wd_in[1030]
  PIN wd_in[1031]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1152.025 0.070 1152.095 ;
    END
  END wd_in[1031]
  PIN wd_in[1032]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1152.165 0.070 1152.235 ;
    END
  END wd_in[1032]
  PIN wd_in[1033]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1152.305 0.070 1152.375 ;
    END
  END wd_in[1033]
  PIN wd_in[1034]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1152.445 0.070 1152.515 ;
    END
  END wd_in[1034]
  PIN wd_in[1035]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1152.585 0.070 1152.655 ;
    END
  END wd_in[1035]
  PIN wd_in[1036]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1152.725 0.070 1152.795 ;
    END
  END wd_in[1036]
  PIN wd_in[1037]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1152.865 0.070 1152.935 ;
    END
  END wd_in[1037]
  PIN wd_in[1038]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.005 0.070 1153.075 ;
    END
  END wd_in[1038]
  PIN wd_in[1039]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.145 0.070 1153.215 ;
    END
  END wd_in[1039]
  PIN wd_in[1040]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.285 0.070 1153.355 ;
    END
  END wd_in[1040]
  PIN wd_in[1041]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.425 0.070 1153.495 ;
    END
  END wd_in[1041]
  PIN wd_in[1042]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.565 0.070 1153.635 ;
    END
  END wd_in[1042]
  PIN wd_in[1043]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.705 0.070 1153.775 ;
    END
  END wd_in[1043]
  PIN wd_in[1044]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.845 0.070 1153.915 ;
    END
  END wd_in[1044]
  PIN wd_in[1045]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1153.985 0.070 1154.055 ;
    END
  END wd_in[1045]
  PIN wd_in[1046]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.125 0.070 1154.195 ;
    END
  END wd_in[1046]
  PIN wd_in[1047]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.265 0.070 1154.335 ;
    END
  END wd_in[1047]
  PIN wd_in[1048]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.405 0.070 1154.475 ;
    END
  END wd_in[1048]
  PIN wd_in[1049]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.545 0.070 1154.615 ;
    END
  END wd_in[1049]
  PIN wd_in[1050]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.685 0.070 1154.755 ;
    END
  END wd_in[1050]
  PIN wd_in[1051]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.825 0.070 1154.895 ;
    END
  END wd_in[1051]
  PIN wd_in[1052]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1154.965 0.070 1155.035 ;
    END
  END wd_in[1052]
  PIN wd_in[1053]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.105 0.070 1155.175 ;
    END
  END wd_in[1053]
  PIN wd_in[1054]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.245 0.070 1155.315 ;
    END
  END wd_in[1054]
  PIN wd_in[1055]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.385 0.070 1155.455 ;
    END
  END wd_in[1055]
  PIN wd_in[1056]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.525 0.070 1155.595 ;
    END
  END wd_in[1056]
  PIN wd_in[1057]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.665 0.070 1155.735 ;
    END
  END wd_in[1057]
  PIN wd_in[1058]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.805 0.070 1155.875 ;
    END
  END wd_in[1058]
  PIN wd_in[1059]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1155.945 0.070 1156.015 ;
    END
  END wd_in[1059]
  PIN wd_in[1060]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1156.085 0.070 1156.155 ;
    END
  END wd_in[1060]
  PIN wd_in[1061]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1156.225 0.070 1156.295 ;
    END
  END wd_in[1061]
  PIN wd_in[1062]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1156.365 0.070 1156.435 ;
    END
  END wd_in[1062]
  PIN wd_in[1063]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1156.505 0.070 1156.575 ;
    END
  END wd_in[1063]
  PIN wd_in[1064]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1156.645 0.070 1156.715 ;
    END
  END wd_in[1064]
  PIN wd_in[1065]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1156.785 0.070 1156.855 ;
    END
  END wd_in[1065]
  PIN wd_in[1066]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1156.925 0.070 1156.995 ;
    END
  END wd_in[1066]
  PIN wd_in[1067]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.065 0.070 1157.135 ;
    END
  END wd_in[1067]
  PIN wd_in[1068]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.205 0.070 1157.275 ;
    END
  END wd_in[1068]
  PIN wd_in[1069]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.345 0.070 1157.415 ;
    END
  END wd_in[1069]
  PIN wd_in[1070]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.485 0.070 1157.555 ;
    END
  END wd_in[1070]
  PIN wd_in[1071]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.625 0.070 1157.695 ;
    END
  END wd_in[1071]
  PIN wd_in[1072]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.765 0.070 1157.835 ;
    END
  END wd_in[1072]
  PIN wd_in[1073]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1157.905 0.070 1157.975 ;
    END
  END wd_in[1073]
  PIN wd_in[1074]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1158.045 0.070 1158.115 ;
    END
  END wd_in[1074]
  PIN wd_in[1075]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1158.185 0.070 1158.255 ;
    END
  END wd_in[1075]
  PIN wd_in[1076]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1158.325 0.070 1158.395 ;
    END
  END wd_in[1076]
  PIN wd_in[1077]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1158.465 0.070 1158.535 ;
    END
  END wd_in[1077]
  PIN wd_in[1078]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1158.605 0.070 1158.675 ;
    END
  END wd_in[1078]
  PIN wd_in[1079]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1158.745 0.070 1158.815 ;
    END
  END wd_in[1079]
  PIN wd_in[1080]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1158.885 0.070 1158.955 ;
    END
  END wd_in[1080]
  PIN wd_in[1081]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1159.025 0.070 1159.095 ;
    END
  END wd_in[1081]
  PIN wd_in[1082]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1159.165 0.070 1159.235 ;
    END
  END wd_in[1082]
  PIN wd_in[1083]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1159.305 0.070 1159.375 ;
    END
  END wd_in[1083]
  PIN wd_in[1084]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1159.445 0.070 1159.515 ;
    END
  END wd_in[1084]
  PIN wd_in[1085]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1159.585 0.070 1159.655 ;
    END
  END wd_in[1085]
  PIN wd_in[1086]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1159.725 0.070 1159.795 ;
    END
  END wd_in[1086]
  PIN wd_in[1087]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1159.865 0.070 1159.935 ;
    END
  END wd_in[1087]
  PIN wd_in[1088]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.005 0.070 1160.075 ;
    END
  END wd_in[1088]
  PIN wd_in[1089]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.145 0.070 1160.215 ;
    END
  END wd_in[1089]
  PIN wd_in[1090]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.285 0.070 1160.355 ;
    END
  END wd_in[1090]
  PIN wd_in[1091]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.425 0.070 1160.495 ;
    END
  END wd_in[1091]
  PIN wd_in[1092]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.565 0.070 1160.635 ;
    END
  END wd_in[1092]
  PIN wd_in[1093]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.705 0.070 1160.775 ;
    END
  END wd_in[1093]
  PIN wd_in[1094]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.845 0.070 1160.915 ;
    END
  END wd_in[1094]
  PIN wd_in[1095]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1160.985 0.070 1161.055 ;
    END
  END wd_in[1095]
  PIN wd_in[1096]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1161.125 0.070 1161.195 ;
    END
  END wd_in[1096]
  PIN wd_in[1097]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1161.265 0.070 1161.335 ;
    END
  END wd_in[1097]
  PIN wd_in[1098]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1161.405 0.070 1161.475 ;
    END
  END wd_in[1098]
  PIN wd_in[1099]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1161.545 0.070 1161.615 ;
    END
  END wd_in[1099]
  PIN wd_in[1100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1161.685 0.070 1161.755 ;
    END
  END wd_in[1100]
  PIN wd_in[1101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1161.825 0.070 1161.895 ;
    END
  END wd_in[1101]
  PIN wd_in[1102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1161.965 0.070 1162.035 ;
    END
  END wd_in[1102]
  PIN wd_in[1103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.105 0.070 1162.175 ;
    END
  END wd_in[1103]
  PIN wd_in[1104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.245 0.070 1162.315 ;
    END
  END wd_in[1104]
  PIN wd_in[1105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.385 0.070 1162.455 ;
    END
  END wd_in[1105]
  PIN wd_in[1106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.525 0.070 1162.595 ;
    END
  END wd_in[1106]
  PIN wd_in[1107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.665 0.070 1162.735 ;
    END
  END wd_in[1107]
  PIN wd_in[1108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.805 0.070 1162.875 ;
    END
  END wd_in[1108]
  PIN wd_in[1109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1162.945 0.070 1163.015 ;
    END
  END wd_in[1109]
  PIN wd_in[1110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1163.085 0.070 1163.155 ;
    END
  END wd_in[1110]
  PIN wd_in[1111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1163.225 0.070 1163.295 ;
    END
  END wd_in[1111]
  PIN wd_in[1112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1163.365 0.070 1163.435 ;
    END
  END wd_in[1112]
  PIN wd_in[1113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1163.505 0.070 1163.575 ;
    END
  END wd_in[1113]
  PIN wd_in[1114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1163.645 0.070 1163.715 ;
    END
  END wd_in[1114]
  PIN wd_in[1115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1163.785 0.070 1163.855 ;
    END
  END wd_in[1115]
  PIN wd_in[1116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1163.925 0.070 1163.995 ;
    END
  END wd_in[1116]
  PIN wd_in[1117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.065 0.070 1164.135 ;
    END
  END wd_in[1117]
  PIN wd_in[1118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.205 0.070 1164.275 ;
    END
  END wd_in[1118]
  PIN wd_in[1119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.345 0.070 1164.415 ;
    END
  END wd_in[1119]
  PIN wd_in[1120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.485 0.070 1164.555 ;
    END
  END wd_in[1120]
  PIN wd_in[1121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.625 0.070 1164.695 ;
    END
  END wd_in[1121]
  PIN wd_in[1122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.765 0.070 1164.835 ;
    END
  END wd_in[1122]
  PIN wd_in[1123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1164.905 0.070 1164.975 ;
    END
  END wd_in[1123]
  PIN wd_in[1124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.045 0.070 1165.115 ;
    END
  END wd_in[1124]
  PIN wd_in[1125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.185 0.070 1165.255 ;
    END
  END wd_in[1125]
  PIN wd_in[1126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.325 0.070 1165.395 ;
    END
  END wd_in[1126]
  PIN wd_in[1127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.465 0.070 1165.535 ;
    END
  END wd_in[1127]
  PIN wd_in[1128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.605 0.070 1165.675 ;
    END
  END wd_in[1128]
  PIN wd_in[1129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.745 0.070 1165.815 ;
    END
  END wd_in[1129]
  PIN wd_in[1130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1165.885 0.070 1165.955 ;
    END
  END wd_in[1130]
  PIN wd_in[1131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1166.025 0.070 1166.095 ;
    END
  END wd_in[1131]
  PIN wd_in[1132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1166.165 0.070 1166.235 ;
    END
  END wd_in[1132]
  PIN wd_in[1133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1166.305 0.070 1166.375 ;
    END
  END wd_in[1133]
  PIN wd_in[1134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1166.445 0.070 1166.515 ;
    END
  END wd_in[1134]
  PIN wd_in[1135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1166.585 0.070 1166.655 ;
    END
  END wd_in[1135]
  PIN wd_in[1136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1166.725 0.070 1166.795 ;
    END
  END wd_in[1136]
  PIN wd_in[1137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1166.865 0.070 1166.935 ;
    END
  END wd_in[1137]
  PIN wd_in[1138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.005 0.070 1167.075 ;
    END
  END wd_in[1138]
  PIN wd_in[1139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.145 0.070 1167.215 ;
    END
  END wd_in[1139]
  PIN wd_in[1140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.285 0.070 1167.355 ;
    END
  END wd_in[1140]
  PIN wd_in[1141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.425 0.070 1167.495 ;
    END
  END wd_in[1141]
  PIN wd_in[1142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.565 0.070 1167.635 ;
    END
  END wd_in[1142]
  PIN wd_in[1143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.705 0.070 1167.775 ;
    END
  END wd_in[1143]
  PIN wd_in[1144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.845 0.070 1167.915 ;
    END
  END wd_in[1144]
  PIN wd_in[1145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1167.985 0.070 1168.055 ;
    END
  END wd_in[1145]
  PIN wd_in[1146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1168.125 0.070 1168.195 ;
    END
  END wd_in[1146]
  PIN wd_in[1147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1168.265 0.070 1168.335 ;
    END
  END wd_in[1147]
  PIN wd_in[1148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1168.405 0.070 1168.475 ;
    END
  END wd_in[1148]
  PIN wd_in[1149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1168.545 0.070 1168.615 ;
    END
  END wd_in[1149]
  PIN wd_in[1150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1168.685 0.070 1168.755 ;
    END
  END wd_in[1150]
  PIN wd_in[1151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1168.825 0.070 1168.895 ;
    END
  END wd_in[1151]
  PIN wd_in[1152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1168.965 0.070 1169.035 ;
    END
  END wd_in[1152]
  PIN wd_in[1153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.105 0.070 1169.175 ;
    END
  END wd_in[1153]
  PIN wd_in[1154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.245 0.070 1169.315 ;
    END
  END wd_in[1154]
  PIN wd_in[1155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.385 0.070 1169.455 ;
    END
  END wd_in[1155]
  PIN wd_in[1156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.525 0.070 1169.595 ;
    END
  END wd_in[1156]
  PIN wd_in[1157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.665 0.070 1169.735 ;
    END
  END wd_in[1157]
  PIN wd_in[1158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.805 0.070 1169.875 ;
    END
  END wd_in[1158]
  PIN wd_in[1159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1169.945 0.070 1170.015 ;
    END
  END wd_in[1159]
  PIN wd_in[1160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1170.085 0.070 1170.155 ;
    END
  END wd_in[1160]
  PIN wd_in[1161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1170.225 0.070 1170.295 ;
    END
  END wd_in[1161]
  PIN wd_in[1162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1170.365 0.070 1170.435 ;
    END
  END wd_in[1162]
  PIN wd_in[1163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1170.505 0.070 1170.575 ;
    END
  END wd_in[1163]
  PIN wd_in[1164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1170.645 0.070 1170.715 ;
    END
  END wd_in[1164]
  PIN wd_in[1165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1170.785 0.070 1170.855 ;
    END
  END wd_in[1165]
  PIN wd_in[1166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1170.925 0.070 1170.995 ;
    END
  END wd_in[1166]
  PIN wd_in[1167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1171.065 0.070 1171.135 ;
    END
  END wd_in[1167]
  PIN wd_in[1168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1171.205 0.070 1171.275 ;
    END
  END wd_in[1168]
  PIN wd_in[1169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1171.345 0.070 1171.415 ;
    END
  END wd_in[1169]
  PIN wd_in[1170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1171.485 0.070 1171.555 ;
    END
  END wd_in[1170]
  PIN wd_in[1171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1171.625 0.070 1171.695 ;
    END
  END wd_in[1171]
  PIN wd_in[1172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1171.765 0.070 1171.835 ;
    END
  END wd_in[1172]
  PIN wd_in[1173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1171.905 0.070 1171.975 ;
    END
  END wd_in[1173]
  PIN wd_in[1174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1172.045 0.070 1172.115 ;
    END
  END wd_in[1174]
  PIN wd_in[1175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1172.185 0.070 1172.255 ;
    END
  END wd_in[1175]
  PIN wd_in[1176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1172.325 0.070 1172.395 ;
    END
  END wd_in[1176]
  PIN wd_in[1177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1172.465 0.070 1172.535 ;
    END
  END wd_in[1177]
  PIN wd_in[1178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1172.605 0.070 1172.675 ;
    END
  END wd_in[1178]
  PIN wd_in[1179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1172.745 0.070 1172.815 ;
    END
  END wd_in[1179]
  PIN wd_in[1180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1172.885 0.070 1172.955 ;
    END
  END wd_in[1180]
  PIN wd_in[1181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1173.025 0.070 1173.095 ;
    END
  END wd_in[1181]
  PIN wd_in[1182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1173.165 0.070 1173.235 ;
    END
  END wd_in[1182]
  PIN wd_in[1183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1173.305 0.070 1173.375 ;
    END
  END wd_in[1183]
  PIN wd_in[1184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1173.445 0.070 1173.515 ;
    END
  END wd_in[1184]
  PIN wd_in[1185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1173.585 0.070 1173.655 ;
    END
  END wd_in[1185]
  PIN wd_in[1186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1173.725 0.070 1173.795 ;
    END
  END wd_in[1186]
  PIN wd_in[1187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1173.865 0.070 1173.935 ;
    END
  END wd_in[1187]
  PIN wd_in[1188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1174.005 0.070 1174.075 ;
    END
  END wd_in[1188]
  PIN wd_in[1189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1174.145 0.070 1174.215 ;
    END
  END wd_in[1189]
  PIN wd_in[1190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1174.285 0.070 1174.355 ;
    END
  END wd_in[1190]
  PIN wd_in[1191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1174.425 0.070 1174.495 ;
    END
  END wd_in[1191]
  PIN wd_in[1192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1174.565 0.070 1174.635 ;
    END
  END wd_in[1192]
  PIN wd_in[1193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1174.705 0.070 1174.775 ;
    END
  END wd_in[1193]
  PIN wd_in[1194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1174.845 0.070 1174.915 ;
    END
  END wd_in[1194]
  PIN wd_in[1195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1174.985 0.070 1175.055 ;
    END
  END wd_in[1195]
  PIN wd_in[1196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1175.125 0.070 1175.195 ;
    END
  END wd_in[1196]
  PIN wd_in[1197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1175.265 0.070 1175.335 ;
    END
  END wd_in[1197]
  PIN wd_in[1198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1175.405 0.070 1175.475 ;
    END
  END wd_in[1198]
  PIN wd_in[1199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1175.545 0.070 1175.615 ;
    END
  END wd_in[1199]
  PIN wd_in[1200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1175.685 0.070 1175.755 ;
    END
  END wd_in[1200]
  PIN wd_in[1201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1175.825 0.070 1175.895 ;
    END
  END wd_in[1201]
  PIN wd_in[1202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1175.965 0.070 1176.035 ;
    END
  END wd_in[1202]
  PIN wd_in[1203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1176.105 0.070 1176.175 ;
    END
  END wd_in[1203]
  PIN wd_in[1204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1176.245 0.070 1176.315 ;
    END
  END wd_in[1204]
  PIN wd_in[1205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1176.385 0.070 1176.455 ;
    END
  END wd_in[1205]
  PIN wd_in[1206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1176.525 0.070 1176.595 ;
    END
  END wd_in[1206]
  PIN wd_in[1207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1176.665 0.070 1176.735 ;
    END
  END wd_in[1207]
  PIN wd_in[1208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1176.805 0.070 1176.875 ;
    END
  END wd_in[1208]
  PIN wd_in[1209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1176.945 0.070 1177.015 ;
    END
  END wd_in[1209]
  PIN wd_in[1210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1177.085 0.070 1177.155 ;
    END
  END wd_in[1210]
  PIN wd_in[1211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1177.225 0.070 1177.295 ;
    END
  END wd_in[1211]
  PIN wd_in[1212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1177.365 0.070 1177.435 ;
    END
  END wd_in[1212]
  PIN wd_in[1213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1177.505 0.070 1177.575 ;
    END
  END wd_in[1213]
  PIN wd_in[1214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1177.645 0.070 1177.715 ;
    END
  END wd_in[1214]
  PIN wd_in[1215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1177.785 0.070 1177.855 ;
    END
  END wd_in[1215]
  PIN wd_in[1216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1177.925 0.070 1177.995 ;
    END
  END wd_in[1216]
  PIN wd_in[1217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1178.065 0.070 1178.135 ;
    END
  END wd_in[1217]
  PIN wd_in[1218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1178.205 0.070 1178.275 ;
    END
  END wd_in[1218]
  PIN wd_in[1219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1178.345 0.070 1178.415 ;
    END
  END wd_in[1219]
  PIN wd_in[1220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1178.485 0.070 1178.555 ;
    END
  END wd_in[1220]
  PIN wd_in[1221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1178.625 0.070 1178.695 ;
    END
  END wd_in[1221]
  PIN wd_in[1222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1178.765 0.070 1178.835 ;
    END
  END wd_in[1222]
  PIN wd_in[1223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1178.905 0.070 1178.975 ;
    END
  END wd_in[1223]
  PIN wd_in[1224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1179.045 0.070 1179.115 ;
    END
  END wd_in[1224]
  PIN wd_in[1225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1179.185 0.070 1179.255 ;
    END
  END wd_in[1225]
  PIN wd_in[1226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1179.325 0.070 1179.395 ;
    END
  END wd_in[1226]
  PIN wd_in[1227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1179.465 0.070 1179.535 ;
    END
  END wd_in[1227]
  PIN wd_in[1228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1179.605 0.070 1179.675 ;
    END
  END wd_in[1228]
  PIN wd_in[1229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1179.745 0.070 1179.815 ;
    END
  END wd_in[1229]
  PIN wd_in[1230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1179.885 0.070 1179.955 ;
    END
  END wd_in[1230]
  PIN wd_in[1231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1180.025 0.070 1180.095 ;
    END
  END wd_in[1231]
  PIN wd_in[1232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1180.165 0.070 1180.235 ;
    END
  END wd_in[1232]
  PIN wd_in[1233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1180.305 0.070 1180.375 ;
    END
  END wd_in[1233]
  PIN wd_in[1234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1180.445 0.070 1180.515 ;
    END
  END wd_in[1234]
  PIN wd_in[1235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1180.585 0.070 1180.655 ;
    END
  END wd_in[1235]
  PIN wd_in[1236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1180.725 0.070 1180.795 ;
    END
  END wd_in[1236]
  PIN wd_in[1237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1180.865 0.070 1180.935 ;
    END
  END wd_in[1237]
  PIN wd_in[1238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1181.005 0.070 1181.075 ;
    END
  END wd_in[1238]
  PIN wd_in[1239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1181.145 0.070 1181.215 ;
    END
  END wd_in[1239]
  PIN wd_in[1240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1181.285 0.070 1181.355 ;
    END
  END wd_in[1240]
  PIN wd_in[1241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1181.425 0.070 1181.495 ;
    END
  END wd_in[1241]
  PIN wd_in[1242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1181.565 0.070 1181.635 ;
    END
  END wd_in[1242]
  PIN wd_in[1243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1181.705 0.070 1181.775 ;
    END
  END wd_in[1243]
  PIN wd_in[1244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1181.845 0.070 1181.915 ;
    END
  END wd_in[1244]
  PIN wd_in[1245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1181.985 0.070 1182.055 ;
    END
  END wd_in[1245]
  PIN wd_in[1246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1182.125 0.070 1182.195 ;
    END
  END wd_in[1246]
  PIN wd_in[1247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1182.265 0.070 1182.335 ;
    END
  END wd_in[1247]
  PIN wd_in[1248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1182.405 0.070 1182.475 ;
    END
  END wd_in[1248]
  PIN wd_in[1249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1182.545 0.070 1182.615 ;
    END
  END wd_in[1249]
  PIN wd_in[1250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1182.685 0.070 1182.755 ;
    END
  END wd_in[1250]
  PIN wd_in[1251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1182.825 0.070 1182.895 ;
    END
  END wd_in[1251]
  PIN wd_in[1252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1182.965 0.070 1183.035 ;
    END
  END wd_in[1252]
  PIN wd_in[1253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1183.105 0.070 1183.175 ;
    END
  END wd_in[1253]
  PIN wd_in[1254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1183.245 0.070 1183.315 ;
    END
  END wd_in[1254]
  PIN wd_in[1255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1183.385 0.070 1183.455 ;
    END
  END wd_in[1255]
  PIN wd_in[1256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1183.525 0.070 1183.595 ;
    END
  END wd_in[1256]
  PIN wd_in[1257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1183.665 0.070 1183.735 ;
    END
  END wd_in[1257]
  PIN wd_in[1258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1183.805 0.070 1183.875 ;
    END
  END wd_in[1258]
  PIN wd_in[1259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1183.945 0.070 1184.015 ;
    END
  END wd_in[1259]
  PIN wd_in[1260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1184.085 0.070 1184.155 ;
    END
  END wd_in[1260]
  PIN wd_in[1261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1184.225 0.070 1184.295 ;
    END
  END wd_in[1261]
  PIN wd_in[1262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1184.365 0.070 1184.435 ;
    END
  END wd_in[1262]
  PIN wd_in[1263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1184.505 0.070 1184.575 ;
    END
  END wd_in[1263]
  PIN wd_in[1264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1184.645 0.070 1184.715 ;
    END
  END wd_in[1264]
  PIN wd_in[1265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1184.785 0.070 1184.855 ;
    END
  END wd_in[1265]
  PIN wd_in[1266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1184.925 0.070 1184.995 ;
    END
  END wd_in[1266]
  PIN wd_in[1267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1185.065 0.070 1185.135 ;
    END
  END wd_in[1267]
  PIN wd_in[1268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1185.205 0.070 1185.275 ;
    END
  END wd_in[1268]
  PIN wd_in[1269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1185.345 0.070 1185.415 ;
    END
  END wd_in[1269]
  PIN wd_in[1270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1185.485 0.070 1185.555 ;
    END
  END wd_in[1270]
  PIN wd_in[1271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1185.625 0.070 1185.695 ;
    END
  END wd_in[1271]
  PIN wd_in[1272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1185.765 0.070 1185.835 ;
    END
  END wd_in[1272]
  PIN wd_in[1273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1185.905 0.070 1185.975 ;
    END
  END wd_in[1273]
  PIN wd_in[1274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1186.045 0.070 1186.115 ;
    END
  END wd_in[1274]
  PIN wd_in[1275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1186.185 0.070 1186.255 ;
    END
  END wd_in[1275]
  PIN wd_in[1276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1186.325 0.070 1186.395 ;
    END
  END wd_in[1276]
  PIN wd_in[1277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1186.465 0.070 1186.535 ;
    END
  END wd_in[1277]
  PIN wd_in[1278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1186.605 0.070 1186.675 ;
    END
  END wd_in[1278]
  PIN wd_in[1279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1186.745 0.070 1186.815 ;
    END
  END wd_in[1279]
  PIN wd_in[1280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1186.885 0.070 1186.955 ;
    END
  END wd_in[1280]
  PIN wd_in[1281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1187.025 0.070 1187.095 ;
    END
  END wd_in[1281]
  PIN wd_in[1282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1187.165 0.070 1187.235 ;
    END
  END wd_in[1282]
  PIN wd_in[1283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1187.305 0.070 1187.375 ;
    END
  END wd_in[1283]
  PIN wd_in[1284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1187.445 0.070 1187.515 ;
    END
  END wd_in[1284]
  PIN wd_in[1285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1187.585 0.070 1187.655 ;
    END
  END wd_in[1285]
  PIN wd_in[1286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1187.725 0.070 1187.795 ;
    END
  END wd_in[1286]
  PIN wd_in[1287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1187.865 0.070 1187.935 ;
    END
  END wd_in[1287]
  PIN wd_in[1288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1188.005 0.070 1188.075 ;
    END
  END wd_in[1288]
  PIN wd_in[1289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1188.145 0.070 1188.215 ;
    END
  END wd_in[1289]
  PIN wd_in[1290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1188.285 0.070 1188.355 ;
    END
  END wd_in[1290]
  PIN wd_in[1291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1188.425 0.070 1188.495 ;
    END
  END wd_in[1291]
  PIN wd_in[1292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1188.565 0.070 1188.635 ;
    END
  END wd_in[1292]
  PIN wd_in[1293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1188.705 0.070 1188.775 ;
    END
  END wd_in[1293]
  PIN wd_in[1294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1188.845 0.070 1188.915 ;
    END
  END wd_in[1294]
  PIN wd_in[1295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1188.985 0.070 1189.055 ;
    END
  END wd_in[1295]
  PIN wd_in[1296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1189.125 0.070 1189.195 ;
    END
  END wd_in[1296]
  PIN wd_in[1297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1189.265 0.070 1189.335 ;
    END
  END wd_in[1297]
  PIN wd_in[1298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1189.405 0.070 1189.475 ;
    END
  END wd_in[1298]
  PIN wd_in[1299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1189.545 0.070 1189.615 ;
    END
  END wd_in[1299]
  PIN wd_in[1300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1189.685 0.070 1189.755 ;
    END
  END wd_in[1300]
  PIN wd_in[1301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1189.825 0.070 1189.895 ;
    END
  END wd_in[1301]
  PIN wd_in[1302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1189.965 0.070 1190.035 ;
    END
  END wd_in[1302]
  PIN wd_in[1303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1190.105 0.070 1190.175 ;
    END
  END wd_in[1303]
  PIN wd_in[1304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1190.245 0.070 1190.315 ;
    END
  END wd_in[1304]
  PIN wd_in[1305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1190.385 0.070 1190.455 ;
    END
  END wd_in[1305]
  PIN wd_in[1306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1190.525 0.070 1190.595 ;
    END
  END wd_in[1306]
  PIN wd_in[1307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1190.665 0.070 1190.735 ;
    END
  END wd_in[1307]
  PIN wd_in[1308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1190.805 0.070 1190.875 ;
    END
  END wd_in[1308]
  PIN wd_in[1309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1190.945 0.070 1191.015 ;
    END
  END wd_in[1309]
  PIN wd_in[1310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1191.085 0.070 1191.155 ;
    END
  END wd_in[1310]
  PIN wd_in[1311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1191.225 0.070 1191.295 ;
    END
  END wd_in[1311]
  PIN wd_in[1312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1191.365 0.070 1191.435 ;
    END
  END wd_in[1312]
  PIN wd_in[1313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1191.505 0.070 1191.575 ;
    END
  END wd_in[1313]
  PIN wd_in[1314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1191.645 0.070 1191.715 ;
    END
  END wd_in[1314]
  PIN wd_in[1315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1191.785 0.070 1191.855 ;
    END
  END wd_in[1315]
  PIN wd_in[1316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1191.925 0.070 1191.995 ;
    END
  END wd_in[1316]
  PIN wd_in[1317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1192.065 0.070 1192.135 ;
    END
  END wd_in[1317]
  PIN wd_in[1318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1192.205 0.070 1192.275 ;
    END
  END wd_in[1318]
  PIN wd_in[1319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1192.345 0.070 1192.415 ;
    END
  END wd_in[1319]
  PIN wd_in[1320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1192.485 0.070 1192.555 ;
    END
  END wd_in[1320]
  PIN wd_in[1321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1192.625 0.070 1192.695 ;
    END
  END wd_in[1321]
  PIN wd_in[1322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1192.765 0.070 1192.835 ;
    END
  END wd_in[1322]
  PIN wd_in[1323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1192.905 0.070 1192.975 ;
    END
  END wd_in[1323]
  PIN wd_in[1324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1193.045 0.070 1193.115 ;
    END
  END wd_in[1324]
  PIN wd_in[1325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1193.185 0.070 1193.255 ;
    END
  END wd_in[1325]
  PIN wd_in[1326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1193.325 0.070 1193.395 ;
    END
  END wd_in[1326]
  PIN wd_in[1327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1193.465 0.070 1193.535 ;
    END
  END wd_in[1327]
  PIN wd_in[1328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1193.605 0.070 1193.675 ;
    END
  END wd_in[1328]
  PIN wd_in[1329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1193.745 0.070 1193.815 ;
    END
  END wd_in[1329]
  PIN wd_in[1330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1193.885 0.070 1193.955 ;
    END
  END wd_in[1330]
  PIN wd_in[1331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1194.025 0.070 1194.095 ;
    END
  END wd_in[1331]
  PIN wd_in[1332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1194.165 0.070 1194.235 ;
    END
  END wd_in[1332]
  PIN wd_in[1333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1194.305 0.070 1194.375 ;
    END
  END wd_in[1333]
  PIN wd_in[1334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1194.445 0.070 1194.515 ;
    END
  END wd_in[1334]
  PIN wd_in[1335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1194.585 0.070 1194.655 ;
    END
  END wd_in[1335]
  PIN wd_in[1336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1194.725 0.070 1194.795 ;
    END
  END wd_in[1336]
  PIN wd_in[1337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1194.865 0.070 1194.935 ;
    END
  END wd_in[1337]
  PIN wd_in[1338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1195.005 0.070 1195.075 ;
    END
  END wd_in[1338]
  PIN wd_in[1339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1195.145 0.070 1195.215 ;
    END
  END wd_in[1339]
  PIN wd_in[1340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1195.285 0.070 1195.355 ;
    END
  END wd_in[1340]
  PIN wd_in[1341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1195.425 0.070 1195.495 ;
    END
  END wd_in[1341]
  PIN wd_in[1342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1195.565 0.070 1195.635 ;
    END
  END wd_in[1342]
  PIN wd_in[1343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1195.705 0.070 1195.775 ;
    END
  END wd_in[1343]
  PIN wd_in[1344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1195.845 0.070 1195.915 ;
    END
  END wd_in[1344]
  PIN wd_in[1345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1195.985 0.070 1196.055 ;
    END
  END wd_in[1345]
  PIN wd_in[1346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1196.125 0.070 1196.195 ;
    END
  END wd_in[1346]
  PIN wd_in[1347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1196.265 0.070 1196.335 ;
    END
  END wd_in[1347]
  PIN wd_in[1348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1196.405 0.070 1196.475 ;
    END
  END wd_in[1348]
  PIN wd_in[1349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1196.545 0.070 1196.615 ;
    END
  END wd_in[1349]
  PIN wd_in[1350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1196.685 0.070 1196.755 ;
    END
  END wd_in[1350]
  PIN wd_in[1351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1196.825 0.070 1196.895 ;
    END
  END wd_in[1351]
  PIN wd_in[1352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1196.965 0.070 1197.035 ;
    END
  END wd_in[1352]
  PIN wd_in[1353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1197.105 0.070 1197.175 ;
    END
  END wd_in[1353]
  PIN wd_in[1354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1197.245 0.070 1197.315 ;
    END
  END wd_in[1354]
  PIN wd_in[1355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1197.385 0.070 1197.455 ;
    END
  END wd_in[1355]
  PIN wd_in[1356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1197.525 0.070 1197.595 ;
    END
  END wd_in[1356]
  PIN wd_in[1357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1197.665 0.070 1197.735 ;
    END
  END wd_in[1357]
  PIN wd_in[1358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1197.805 0.070 1197.875 ;
    END
  END wd_in[1358]
  PIN wd_in[1359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1197.945 0.070 1198.015 ;
    END
  END wd_in[1359]
  PIN wd_in[1360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1198.085 0.070 1198.155 ;
    END
  END wd_in[1360]
  PIN wd_in[1361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1198.225 0.070 1198.295 ;
    END
  END wd_in[1361]
  PIN wd_in[1362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1198.365 0.070 1198.435 ;
    END
  END wd_in[1362]
  PIN wd_in[1363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1198.505 0.070 1198.575 ;
    END
  END wd_in[1363]
  PIN wd_in[1364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1198.645 0.070 1198.715 ;
    END
  END wd_in[1364]
  PIN wd_in[1365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1198.785 0.070 1198.855 ;
    END
  END wd_in[1365]
  PIN wd_in[1366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1198.925 0.070 1198.995 ;
    END
  END wd_in[1366]
  PIN wd_in[1367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1199.065 0.070 1199.135 ;
    END
  END wd_in[1367]
  PIN wd_in[1368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1199.205 0.070 1199.275 ;
    END
  END wd_in[1368]
  PIN wd_in[1369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1199.345 0.070 1199.415 ;
    END
  END wd_in[1369]
  PIN wd_in[1370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1199.485 0.070 1199.555 ;
    END
  END wd_in[1370]
  PIN wd_in[1371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1199.625 0.070 1199.695 ;
    END
  END wd_in[1371]
  PIN wd_in[1372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1199.765 0.070 1199.835 ;
    END
  END wd_in[1372]
  PIN wd_in[1373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1199.905 0.070 1199.975 ;
    END
  END wd_in[1373]
  PIN wd_in[1374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1200.045 0.070 1200.115 ;
    END
  END wd_in[1374]
  PIN wd_in[1375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1200.185 0.070 1200.255 ;
    END
  END wd_in[1375]
  PIN wd_in[1376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1200.325 0.070 1200.395 ;
    END
  END wd_in[1376]
  PIN wd_in[1377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1200.465 0.070 1200.535 ;
    END
  END wd_in[1377]
  PIN wd_in[1378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1200.605 0.070 1200.675 ;
    END
  END wd_in[1378]
  PIN wd_in[1379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1200.745 0.070 1200.815 ;
    END
  END wd_in[1379]
  PIN wd_in[1380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1200.885 0.070 1200.955 ;
    END
  END wd_in[1380]
  PIN wd_in[1381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1201.025 0.070 1201.095 ;
    END
  END wd_in[1381]
  PIN wd_in[1382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1201.165 0.070 1201.235 ;
    END
  END wd_in[1382]
  PIN wd_in[1383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1201.305 0.070 1201.375 ;
    END
  END wd_in[1383]
  PIN wd_in[1384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1201.445 0.070 1201.515 ;
    END
  END wd_in[1384]
  PIN wd_in[1385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1201.585 0.070 1201.655 ;
    END
  END wd_in[1385]
  PIN wd_in[1386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1201.725 0.070 1201.795 ;
    END
  END wd_in[1386]
  PIN wd_in[1387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1201.865 0.070 1201.935 ;
    END
  END wd_in[1387]
  PIN wd_in[1388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1202.005 0.070 1202.075 ;
    END
  END wd_in[1388]
  PIN wd_in[1389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1202.145 0.070 1202.215 ;
    END
  END wd_in[1389]
  PIN wd_in[1390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1202.285 0.070 1202.355 ;
    END
  END wd_in[1390]
  PIN wd_in[1391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1202.425 0.070 1202.495 ;
    END
  END wd_in[1391]
  PIN wd_in[1392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1202.565 0.070 1202.635 ;
    END
  END wd_in[1392]
  PIN wd_in[1393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1202.705 0.070 1202.775 ;
    END
  END wd_in[1393]
  PIN wd_in[1394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1202.845 0.070 1202.915 ;
    END
  END wd_in[1394]
  PIN wd_in[1395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1202.985 0.070 1203.055 ;
    END
  END wd_in[1395]
  PIN wd_in[1396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1203.125 0.070 1203.195 ;
    END
  END wd_in[1396]
  PIN wd_in[1397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1203.265 0.070 1203.335 ;
    END
  END wd_in[1397]
  PIN wd_in[1398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1203.405 0.070 1203.475 ;
    END
  END wd_in[1398]
  PIN wd_in[1399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1203.545 0.070 1203.615 ;
    END
  END wd_in[1399]
  PIN wd_in[1400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1203.685 0.070 1203.755 ;
    END
  END wd_in[1400]
  PIN wd_in[1401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1203.825 0.070 1203.895 ;
    END
  END wd_in[1401]
  PIN wd_in[1402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1203.965 0.070 1204.035 ;
    END
  END wd_in[1402]
  PIN wd_in[1403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1204.105 0.070 1204.175 ;
    END
  END wd_in[1403]
  PIN wd_in[1404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1204.245 0.070 1204.315 ;
    END
  END wd_in[1404]
  PIN wd_in[1405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1204.385 0.070 1204.455 ;
    END
  END wd_in[1405]
  PIN wd_in[1406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1204.525 0.070 1204.595 ;
    END
  END wd_in[1406]
  PIN wd_in[1407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1204.665 0.070 1204.735 ;
    END
  END wd_in[1407]
  PIN wd_in[1408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1204.805 0.070 1204.875 ;
    END
  END wd_in[1408]
  PIN wd_in[1409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1204.945 0.070 1205.015 ;
    END
  END wd_in[1409]
  PIN wd_in[1410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1205.085 0.070 1205.155 ;
    END
  END wd_in[1410]
  PIN wd_in[1411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1205.225 0.070 1205.295 ;
    END
  END wd_in[1411]
  PIN wd_in[1412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1205.365 0.070 1205.435 ;
    END
  END wd_in[1412]
  PIN wd_in[1413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1205.505 0.070 1205.575 ;
    END
  END wd_in[1413]
  PIN wd_in[1414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1205.645 0.070 1205.715 ;
    END
  END wd_in[1414]
  PIN wd_in[1415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1205.785 0.070 1205.855 ;
    END
  END wd_in[1415]
  PIN wd_in[1416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1205.925 0.070 1205.995 ;
    END
  END wd_in[1416]
  PIN wd_in[1417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1206.065 0.070 1206.135 ;
    END
  END wd_in[1417]
  PIN wd_in[1418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1206.205 0.070 1206.275 ;
    END
  END wd_in[1418]
  PIN wd_in[1419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1206.345 0.070 1206.415 ;
    END
  END wd_in[1419]
  PIN wd_in[1420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1206.485 0.070 1206.555 ;
    END
  END wd_in[1420]
  PIN wd_in[1421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1206.625 0.070 1206.695 ;
    END
  END wd_in[1421]
  PIN wd_in[1422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1206.765 0.070 1206.835 ;
    END
  END wd_in[1422]
  PIN wd_in[1423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1206.905 0.070 1206.975 ;
    END
  END wd_in[1423]
  PIN wd_in[1424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1207.045 0.070 1207.115 ;
    END
  END wd_in[1424]
  PIN wd_in[1425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1207.185 0.070 1207.255 ;
    END
  END wd_in[1425]
  PIN wd_in[1426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1207.325 0.070 1207.395 ;
    END
  END wd_in[1426]
  PIN wd_in[1427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1207.465 0.070 1207.535 ;
    END
  END wd_in[1427]
  PIN wd_in[1428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1207.605 0.070 1207.675 ;
    END
  END wd_in[1428]
  PIN wd_in[1429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1207.745 0.070 1207.815 ;
    END
  END wd_in[1429]
  PIN wd_in[1430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1207.885 0.070 1207.955 ;
    END
  END wd_in[1430]
  PIN wd_in[1431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1208.025 0.070 1208.095 ;
    END
  END wd_in[1431]
  PIN wd_in[1432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1208.165 0.070 1208.235 ;
    END
  END wd_in[1432]
  PIN wd_in[1433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1208.305 0.070 1208.375 ;
    END
  END wd_in[1433]
  PIN wd_in[1434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1208.445 0.070 1208.515 ;
    END
  END wd_in[1434]
  PIN wd_in[1435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1208.585 0.070 1208.655 ;
    END
  END wd_in[1435]
  PIN wd_in[1436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1208.725 0.070 1208.795 ;
    END
  END wd_in[1436]
  PIN wd_in[1437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1208.865 0.070 1208.935 ;
    END
  END wd_in[1437]
  PIN wd_in[1438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1209.005 0.070 1209.075 ;
    END
  END wd_in[1438]
  PIN wd_in[1439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1209.145 0.070 1209.215 ;
    END
  END wd_in[1439]
  PIN wd_in[1440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1209.285 0.070 1209.355 ;
    END
  END wd_in[1440]
  PIN wd_in[1441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1209.425 0.070 1209.495 ;
    END
  END wd_in[1441]
  PIN wd_in[1442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1209.565 0.070 1209.635 ;
    END
  END wd_in[1442]
  PIN wd_in[1443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1209.705 0.070 1209.775 ;
    END
  END wd_in[1443]
  PIN wd_in[1444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1209.845 0.070 1209.915 ;
    END
  END wd_in[1444]
  PIN wd_in[1445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1209.985 0.070 1210.055 ;
    END
  END wd_in[1445]
  PIN wd_in[1446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1210.125 0.070 1210.195 ;
    END
  END wd_in[1446]
  PIN wd_in[1447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1210.265 0.070 1210.335 ;
    END
  END wd_in[1447]
  PIN wd_in[1448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1210.405 0.070 1210.475 ;
    END
  END wd_in[1448]
  PIN wd_in[1449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1210.545 0.070 1210.615 ;
    END
  END wd_in[1449]
  PIN wd_in[1450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1210.685 0.070 1210.755 ;
    END
  END wd_in[1450]
  PIN wd_in[1451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1210.825 0.070 1210.895 ;
    END
  END wd_in[1451]
  PIN wd_in[1452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1210.965 0.070 1211.035 ;
    END
  END wd_in[1452]
  PIN wd_in[1453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1211.105 0.070 1211.175 ;
    END
  END wd_in[1453]
  PIN wd_in[1454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1211.245 0.070 1211.315 ;
    END
  END wd_in[1454]
  PIN wd_in[1455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1211.385 0.070 1211.455 ;
    END
  END wd_in[1455]
  PIN wd_in[1456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1211.525 0.070 1211.595 ;
    END
  END wd_in[1456]
  PIN wd_in[1457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1211.665 0.070 1211.735 ;
    END
  END wd_in[1457]
  PIN wd_in[1458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1211.805 0.070 1211.875 ;
    END
  END wd_in[1458]
  PIN wd_in[1459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1211.945 0.070 1212.015 ;
    END
  END wd_in[1459]
  PIN wd_in[1460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1212.085 0.070 1212.155 ;
    END
  END wd_in[1460]
  PIN wd_in[1461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1212.225 0.070 1212.295 ;
    END
  END wd_in[1461]
  PIN wd_in[1462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1212.365 0.070 1212.435 ;
    END
  END wd_in[1462]
  PIN wd_in[1463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1212.505 0.070 1212.575 ;
    END
  END wd_in[1463]
  PIN wd_in[1464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1212.645 0.070 1212.715 ;
    END
  END wd_in[1464]
  PIN wd_in[1465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1212.785 0.070 1212.855 ;
    END
  END wd_in[1465]
  PIN wd_in[1466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1212.925 0.070 1212.995 ;
    END
  END wd_in[1466]
  PIN wd_in[1467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1213.065 0.070 1213.135 ;
    END
  END wd_in[1467]
  PIN wd_in[1468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1213.205 0.070 1213.275 ;
    END
  END wd_in[1468]
  PIN wd_in[1469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1213.345 0.070 1213.415 ;
    END
  END wd_in[1469]
  PIN wd_in[1470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1213.485 0.070 1213.555 ;
    END
  END wd_in[1470]
  PIN wd_in[1471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1213.625 0.070 1213.695 ;
    END
  END wd_in[1471]
  PIN wd_in[1472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1213.765 0.070 1213.835 ;
    END
  END wd_in[1472]
  PIN wd_in[1473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1213.905 0.070 1213.975 ;
    END
  END wd_in[1473]
  PIN wd_in[1474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1214.045 0.070 1214.115 ;
    END
  END wd_in[1474]
  PIN wd_in[1475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1214.185 0.070 1214.255 ;
    END
  END wd_in[1475]
  PIN wd_in[1476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1214.325 0.070 1214.395 ;
    END
  END wd_in[1476]
  PIN wd_in[1477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1214.465 0.070 1214.535 ;
    END
  END wd_in[1477]
  PIN wd_in[1478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1214.605 0.070 1214.675 ;
    END
  END wd_in[1478]
  PIN wd_in[1479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1214.745 0.070 1214.815 ;
    END
  END wd_in[1479]
  PIN wd_in[1480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1214.885 0.070 1214.955 ;
    END
  END wd_in[1480]
  PIN wd_in[1481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1215.025 0.070 1215.095 ;
    END
  END wd_in[1481]
  PIN wd_in[1482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1215.165 0.070 1215.235 ;
    END
  END wd_in[1482]
  PIN wd_in[1483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1215.305 0.070 1215.375 ;
    END
  END wd_in[1483]
  PIN wd_in[1484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1215.445 0.070 1215.515 ;
    END
  END wd_in[1484]
  PIN wd_in[1485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1215.585 0.070 1215.655 ;
    END
  END wd_in[1485]
  PIN wd_in[1486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1215.725 0.070 1215.795 ;
    END
  END wd_in[1486]
  PIN wd_in[1487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1215.865 0.070 1215.935 ;
    END
  END wd_in[1487]
  PIN wd_in[1488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1216.005 0.070 1216.075 ;
    END
  END wd_in[1488]
  PIN wd_in[1489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1216.145 0.070 1216.215 ;
    END
  END wd_in[1489]
  PIN wd_in[1490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1216.285 0.070 1216.355 ;
    END
  END wd_in[1490]
  PIN wd_in[1491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1216.425 0.070 1216.495 ;
    END
  END wd_in[1491]
  PIN wd_in[1492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1216.565 0.070 1216.635 ;
    END
  END wd_in[1492]
  PIN wd_in[1493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1216.705 0.070 1216.775 ;
    END
  END wd_in[1493]
  PIN wd_in[1494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1216.845 0.070 1216.915 ;
    END
  END wd_in[1494]
  PIN wd_in[1495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1216.985 0.070 1217.055 ;
    END
  END wd_in[1495]
  PIN wd_in[1496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1217.125 0.070 1217.195 ;
    END
  END wd_in[1496]
  PIN wd_in[1497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1217.265 0.070 1217.335 ;
    END
  END wd_in[1497]
  PIN wd_in[1498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1217.405 0.070 1217.475 ;
    END
  END wd_in[1498]
  PIN wd_in[1499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1217.545 0.070 1217.615 ;
    END
  END wd_in[1499]
  PIN wd_in[1500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1217.685 0.070 1217.755 ;
    END
  END wd_in[1500]
  PIN wd_in[1501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1217.825 0.070 1217.895 ;
    END
  END wd_in[1501]
  PIN wd_in[1502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1217.965 0.070 1218.035 ;
    END
  END wd_in[1502]
  PIN wd_in[1503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.105 0.070 1218.175 ;
    END
  END wd_in[1503]
  PIN wd_in[1504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.245 0.070 1218.315 ;
    END
  END wd_in[1504]
  PIN wd_in[1505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.385 0.070 1218.455 ;
    END
  END wd_in[1505]
  PIN wd_in[1506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.525 0.070 1218.595 ;
    END
  END wd_in[1506]
  PIN wd_in[1507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.665 0.070 1218.735 ;
    END
  END wd_in[1507]
  PIN wd_in[1508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.805 0.070 1218.875 ;
    END
  END wd_in[1508]
  PIN wd_in[1509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1218.945 0.070 1219.015 ;
    END
  END wd_in[1509]
  PIN wd_in[1510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.085 0.070 1219.155 ;
    END
  END wd_in[1510]
  PIN wd_in[1511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.225 0.070 1219.295 ;
    END
  END wd_in[1511]
  PIN wd_in[1512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.365 0.070 1219.435 ;
    END
  END wd_in[1512]
  PIN wd_in[1513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.505 0.070 1219.575 ;
    END
  END wd_in[1513]
  PIN wd_in[1514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.645 0.070 1219.715 ;
    END
  END wd_in[1514]
  PIN wd_in[1515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.785 0.070 1219.855 ;
    END
  END wd_in[1515]
  PIN wd_in[1516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1219.925 0.070 1219.995 ;
    END
  END wd_in[1516]
  PIN wd_in[1517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1220.065 0.070 1220.135 ;
    END
  END wd_in[1517]
  PIN wd_in[1518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1220.205 0.070 1220.275 ;
    END
  END wd_in[1518]
  PIN wd_in[1519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1220.345 0.070 1220.415 ;
    END
  END wd_in[1519]
  PIN wd_in[1520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1220.485 0.070 1220.555 ;
    END
  END wd_in[1520]
  PIN wd_in[1521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1220.625 0.070 1220.695 ;
    END
  END wd_in[1521]
  PIN wd_in[1522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1220.765 0.070 1220.835 ;
    END
  END wd_in[1522]
  PIN wd_in[1523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1220.905 0.070 1220.975 ;
    END
  END wd_in[1523]
  PIN wd_in[1524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1221.045 0.070 1221.115 ;
    END
  END wd_in[1524]
  PIN wd_in[1525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1221.185 0.070 1221.255 ;
    END
  END wd_in[1525]
  PIN wd_in[1526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1221.325 0.070 1221.395 ;
    END
  END wd_in[1526]
  PIN wd_in[1527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1221.465 0.070 1221.535 ;
    END
  END wd_in[1527]
  PIN wd_in[1528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1221.605 0.070 1221.675 ;
    END
  END wd_in[1528]
  PIN wd_in[1529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1221.745 0.070 1221.815 ;
    END
  END wd_in[1529]
  PIN wd_in[1530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1221.885 0.070 1221.955 ;
    END
  END wd_in[1530]
  PIN wd_in[1531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.025 0.070 1222.095 ;
    END
  END wd_in[1531]
  PIN wd_in[1532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.165 0.070 1222.235 ;
    END
  END wd_in[1532]
  PIN wd_in[1533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.305 0.070 1222.375 ;
    END
  END wd_in[1533]
  PIN wd_in[1534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.445 0.070 1222.515 ;
    END
  END wd_in[1534]
  PIN wd_in[1535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.585 0.070 1222.655 ;
    END
  END wd_in[1535]
  PIN wd_in[1536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.725 0.070 1222.795 ;
    END
  END wd_in[1536]
  PIN wd_in[1537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1222.865 0.070 1222.935 ;
    END
  END wd_in[1537]
  PIN wd_in[1538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.005 0.070 1223.075 ;
    END
  END wd_in[1538]
  PIN wd_in[1539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.145 0.070 1223.215 ;
    END
  END wd_in[1539]
  PIN wd_in[1540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.285 0.070 1223.355 ;
    END
  END wd_in[1540]
  PIN wd_in[1541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.425 0.070 1223.495 ;
    END
  END wd_in[1541]
  PIN wd_in[1542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.565 0.070 1223.635 ;
    END
  END wd_in[1542]
  PIN wd_in[1543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.705 0.070 1223.775 ;
    END
  END wd_in[1543]
  PIN wd_in[1544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.845 0.070 1223.915 ;
    END
  END wd_in[1544]
  PIN wd_in[1545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1223.985 0.070 1224.055 ;
    END
  END wd_in[1545]
  PIN wd_in[1546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.125 0.070 1224.195 ;
    END
  END wd_in[1546]
  PIN wd_in[1547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.265 0.070 1224.335 ;
    END
  END wd_in[1547]
  PIN wd_in[1548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.405 0.070 1224.475 ;
    END
  END wd_in[1548]
  PIN wd_in[1549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.545 0.070 1224.615 ;
    END
  END wd_in[1549]
  PIN wd_in[1550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.685 0.070 1224.755 ;
    END
  END wd_in[1550]
  PIN wd_in[1551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.825 0.070 1224.895 ;
    END
  END wd_in[1551]
  PIN wd_in[1552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1224.965 0.070 1225.035 ;
    END
  END wd_in[1552]
  PIN wd_in[1553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1225.105 0.070 1225.175 ;
    END
  END wd_in[1553]
  PIN wd_in[1554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1225.245 0.070 1225.315 ;
    END
  END wd_in[1554]
  PIN wd_in[1555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1225.385 0.070 1225.455 ;
    END
  END wd_in[1555]
  PIN wd_in[1556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1225.525 0.070 1225.595 ;
    END
  END wd_in[1556]
  PIN wd_in[1557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1225.665 0.070 1225.735 ;
    END
  END wd_in[1557]
  PIN wd_in[1558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1225.805 0.070 1225.875 ;
    END
  END wd_in[1558]
  PIN wd_in[1559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1225.945 0.070 1226.015 ;
    END
  END wd_in[1559]
  PIN wd_in[1560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1226.085 0.070 1226.155 ;
    END
  END wd_in[1560]
  PIN wd_in[1561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1226.225 0.070 1226.295 ;
    END
  END wd_in[1561]
  PIN wd_in[1562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1226.365 0.070 1226.435 ;
    END
  END wd_in[1562]
  PIN wd_in[1563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1226.505 0.070 1226.575 ;
    END
  END wd_in[1563]
  PIN wd_in[1564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1226.645 0.070 1226.715 ;
    END
  END wd_in[1564]
  PIN wd_in[1565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1226.785 0.070 1226.855 ;
    END
  END wd_in[1565]
  PIN wd_in[1566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1226.925 0.070 1226.995 ;
    END
  END wd_in[1566]
  PIN wd_in[1567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1227.065 0.070 1227.135 ;
    END
  END wd_in[1567]
  PIN wd_in[1568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1227.205 0.070 1227.275 ;
    END
  END wd_in[1568]
  PIN wd_in[1569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1227.345 0.070 1227.415 ;
    END
  END wd_in[1569]
  PIN wd_in[1570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1227.485 0.070 1227.555 ;
    END
  END wd_in[1570]
  PIN wd_in[1571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1227.625 0.070 1227.695 ;
    END
  END wd_in[1571]
  PIN wd_in[1572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1227.765 0.070 1227.835 ;
    END
  END wd_in[1572]
  PIN wd_in[1573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1227.905 0.070 1227.975 ;
    END
  END wd_in[1573]
  PIN wd_in[1574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1228.045 0.070 1228.115 ;
    END
  END wd_in[1574]
  PIN wd_in[1575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1228.185 0.070 1228.255 ;
    END
  END wd_in[1575]
  PIN wd_in[1576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1228.325 0.070 1228.395 ;
    END
  END wd_in[1576]
  PIN wd_in[1577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1228.465 0.070 1228.535 ;
    END
  END wd_in[1577]
  PIN wd_in[1578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1228.605 0.070 1228.675 ;
    END
  END wd_in[1578]
  PIN wd_in[1579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1228.745 0.070 1228.815 ;
    END
  END wd_in[1579]
  PIN wd_in[1580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1228.885 0.070 1228.955 ;
    END
  END wd_in[1580]
  PIN wd_in[1581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1229.025 0.070 1229.095 ;
    END
  END wd_in[1581]
  PIN wd_in[1582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1229.165 0.070 1229.235 ;
    END
  END wd_in[1582]
  PIN wd_in[1583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1229.305 0.070 1229.375 ;
    END
  END wd_in[1583]
  PIN wd_in[1584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1229.445 0.070 1229.515 ;
    END
  END wd_in[1584]
  PIN wd_in[1585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1229.585 0.070 1229.655 ;
    END
  END wd_in[1585]
  PIN wd_in[1586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1229.725 0.070 1229.795 ;
    END
  END wd_in[1586]
  PIN wd_in[1587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1229.865 0.070 1229.935 ;
    END
  END wd_in[1587]
  PIN wd_in[1588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1230.005 0.070 1230.075 ;
    END
  END wd_in[1588]
  PIN wd_in[1589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1230.145 0.070 1230.215 ;
    END
  END wd_in[1589]
  PIN wd_in[1590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1230.285 0.070 1230.355 ;
    END
  END wd_in[1590]
  PIN wd_in[1591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1230.425 0.070 1230.495 ;
    END
  END wd_in[1591]
  PIN wd_in[1592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1230.565 0.070 1230.635 ;
    END
  END wd_in[1592]
  PIN wd_in[1593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1230.705 0.070 1230.775 ;
    END
  END wd_in[1593]
  PIN wd_in[1594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1230.845 0.070 1230.915 ;
    END
  END wd_in[1594]
  PIN wd_in[1595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1230.985 0.070 1231.055 ;
    END
  END wd_in[1595]
  PIN wd_in[1596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1231.125 0.070 1231.195 ;
    END
  END wd_in[1596]
  PIN wd_in[1597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1231.265 0.070 1231.335 ;
    END
  END wd_in[1597]
  PIN wd_in[1598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1231.405 0.070 1231.475 ;
    END
  END wd_in[1598]
  PIN wd_in[1599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1231.545 0.070 1231.615 ;
    END
  END wd_in[1599]
  PIN wd_in[1600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1231.685 0.070 1231.755 ;
    END
  END wd_in[1600]
  PIN wd_in[1601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1231.825 0.070 1231.895 ;
    END
  END wd_in[1601]
  PIN wd_in[1602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1231.965 0.070 1232.035 ;
    END
  END wd_in[1602]
  PIN wd_in[1603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1232.105 0.070 1232.175 ;
    END
  END wd_in[1603]
  PIN wd_in[1604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1232.245 0.070 1232.315 ;
    END
  END wd_in[1604]
  PIN wd_in[1605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1232.385 0.070 1232.455 ;
    END
  END wd_in[1605]
  PIN wd_in[1606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1232.525 0.070 1232.595 ;
    END
  END wd_in[1606]
  PIN wd_in[1607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1232.665 0.070 1232.735 ;
    END
  END wd_in[1607]
  PIN wd_in[1608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1232.805 0.070 1232.875 ;
    END
  END wd_in[1608]
  PIN wd_in[1609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1232.945 0.070 1233.015 ;
    END
  END wd_in[1609]
  PIN wd_in[1610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1233.085 0.070 1233.155 ;
    END
  END wd_in[1610]
  PIN wd_in[1611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1233.225 0.070 1233.295 ;
    END
  END wd_in[1611]
  PIN wd_in[1612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1233.365 0.070 1233.435 ;
    END
  END wd_in[1612]
  PIN wd_in[1613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1233.505 0.070 1233.575 ;
    END
  END wd_in[1613]
  PIN wd_in[1614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1233.645 0.070 1233.715 ;
    END
  END wd_in[1614]
  PIN wd_in[1615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1233.785 0.070 1233.855 ;
    END
  END wd_in[1615]
  PIN wd_in[1616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1233.925 0.070 1233.995 ;
    END
  END wd_in[1616]
  PIN wd_in[1617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1234.065 0.070 1234.135 ;
    END
  END wd_in[1617]
  PIN wd_in[1618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1234.205 0.070 1234.275 ;
    END
  END wd_in[1618]
  PIN wd_in[1619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1234.345 0.070 1234.415 ;
    END
  END wd_in[1619]
  PIN wd_in[1620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1234.485 0.070 1234.555 ;
    END
  END wd_in[1620]
  PIN wd_in[1621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1234.625 0.070 1234.695 ;
    END
  END wd_in[1621]
  PIN wd_in[1622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1234.765 0.070 1234.835 ;
    END
  END wd_in[1622]
  PIN wd_in[1623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1234.905 0.070 1234.975 ;
    END
  END wd_in[1623]
  PIN wd_in[1624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1235.045 0.070 1235.115 ;
    END
  END wd_in[1624]
  PIN wd_in[1625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1235.185 0.070 1235.255 ;
    END
  END wd_in[1625]
  PIN wd_in[1626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1235.325 0.070 1235.395 ;
    END
  END wd_in[1626]
  PIN wd_in[1627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1235.465 0.070 1235.535 ;
    END
  END wd_in[1627]
  PIN wd_in[1628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1235.605 0.070 1235.675 ;
    END
  END wd_in[1628]
  PIN wd_in[1629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1235.745 0.070 1235.815 ;
    END
  END wd_in[1629]
  PIN wd_in[1630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1235.885 0.070 1235.955 ;
    END
  END wd_in[1630]
  PIN wd_in[1631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1236.025 0.070 1236.095 ;
    END
  END wd_in[1631]
  PIN wd_in[1632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1236.165 0.070 1236.235 ;
    END
  END wd_in[1632]
  PIN wd_in[1633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1236.305 0.070 1236.375 ;
    END
  END wd_in[1633]
  PIN wd_in[1634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1236.445 0.070 1236.515 ;
    END
  END wd_in[1634]
  PIN wd_in[1635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1236.585 0.070 1236.655 ;
    END
  END wd_in[1635]
  PIN wd_in[1636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1236.725 0.070 1236.795 ;
    END
  END wd_in[1636]
  PIN wd_in[1637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1236.865 0.070 1236.935 ;
    END
  END wd_in[1637]
  PIN wd_in[1638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1237.005 0.070 1237.075 ;
    END
  END wd_in[1638]
  PIN wd_in[1639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1237.145 0.070 1237.215 ;
    END
  END wd_in[1639]
  PIN wd_in[1640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1237.285 0.070 1237.355 ;
    END
  END wd_in[1640]
  PIN wd_in[1641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1237.425 0.070 1237.495 ;
    END
  END wd_in[1641]
  PIN wd_in[1642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1237.565 0.070 1237.635 ;
    END
  END wd_in[1642]
  PIN wd_in[1643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1237.705 0.070 1237.775 ;
    END
  END wd_in[1643]
  PIN wd_in[1644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1237.845 0.070 1237.915 ;
    END
  END wd_in[1644]
  PIN wd_in[1645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1237.985 0.070 1238.055 ;
    END
  END wd_in[1645]
  PIN wd_in[1646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1238.125 0.070 1238.195 ;
    END
  END wd_in[1646]
  PIN wd_in[1647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1238.265 0.070 1238.335 ;
    END
  END wd_in[1647]
  PIN wd_in[1648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1238.405 0.070 1238.475 ;
    END
  END wd_in[1648]
  PIN wd_in[1649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1238.545 0.070 1238.615 ;
    END
  END wd_in[1649]
  PIN wd_in[1650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1238.685 0.070 1238.755 ;
    END
  END wd_in[1650]
  PIN wd_in[1651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1238.825 0.070 1238.895 ;
    END
  END wd_in[1651]
  PIN wd_in[1652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1238.965 0.070 1239.035 ;
    END
  END wd_in[1652]
  PIN wd_in[1653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1239.105 0.070 1239.175 ;
    END
  END wd_in[1653]
  PIN wd_in[1654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1239.245 0.070 1239.315 ;
    END
  END wd_in[1654]
  PIN wd_in[1655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1239.385 0.070 1239.455 ;
    END
  END wd_in[1655]
  PIN wd_in[1656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1239.525 0.070 1239.595 ;
    END
  END wd_in[1656]
  PIN wd_in[1657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1239.665 0.070 1239.735 ;
    END
  END wd_in[1657]
  PIN wd_in[1658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1239.805 0.070 1239.875 ;
    END
  END wd_in[1658]
  PIN wd_in[1659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1239.945 0.070 1240.015 ;
    END
  END wd_in[1659]
  PIN wd_in[1660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1240.085 0.070 1240.155 ;
    END
  END wd_in[1660]
  PIN wd_in[1661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1240.225 0.070 1240.295 ;
    END
  END wd_in[1661]
  PIN wd_in[1662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1240.365 0.070 1240.435 ;
    END
  END wd_in[1662]
  PIN wd_in[1663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1240.505 0.070 1240.575 ;
    END
  END wd_in[1663]
  PIN wd_in[1664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1240.645 0.070 1240.715 ;
    END
  END wd_in[1664]
  PIN wd_in[1665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1240.785 0.070 1240.855 ;
    END
  END wd_in[1665]
  PIN wd_in[1666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1240.925 0.070 1240.995 ;
    END
  END wd_in[1666]
  PIN wd_in[1667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1241.065 0.070 1241.135 ;
    END
  END wd_in[1667]
  PIN wd_in[1668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1241.205 0.070 1241.275 ;
    END
  END wd_in[1668]
  PIN wd_in[1669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1241.345 0.070 1241.415 ;
    END
  END wd_in[1669]
  PIN wd_in[1670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1241.485 0.070 1241.555 ;
    END
  END wd_in[1670]
  PIN wd_in[1671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1241.625 0.070 1241.695 ;
    END
  END wd_in[1671]
  PIN wd_in[1672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1241.765 0.070 1241.835 ;
    END
  END wd_in[1672]
  PIN wd_in[1673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1241.905 0.070 1241.975 ;
    END
  END wd_in[1673]
  PIN wd_in[1674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1242.045 0.070 1242.115 ;
    END
  END wd_in[1674]
  PIN wd_in[1675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1242.185 0.070 1242.255 ;
    END
  END wd_in[1675]
  PIN wd_in[1676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1242.325 0.070 1242.395 ;
    END
  END wd_in[1676]
  PIN wd_in[1677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1242.465 0.070 1242.535 ;
    END
  END wd_in[1677]
  PIN wd_in[1678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1242.605 0.070 1242.675 ;
    END
  END wd_in[1678]
  PIN wd_in[1679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1242.745 0.070 1242.815 ;
    END
  END wd_in[1679]
  PIN wd_in[1680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1242.885 0.070 1242.955 ;
    END
  END wd_in[1680]
  PIN wd_in[1681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1243.025 0.070 1243.095 ;
    END
  END wd_in[1681]
  PIN wd_in[1682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1243.165 0.070 1243.235 ;
    END
  END wd_in[1682]
  PIN wd_in[1683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1243.305 0.070 1243.375 ;
    END
  END wd_in[1683]
  PIN wd_in[1684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1243.445 0.070 1243.515 ;
    END
  END wd_in[1684]
  PIN wd_in[1685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1243.585 0.070 1243.655 ;
    END
  END wd_in[1685]
  PIN wd_in[1686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1243.725 0.070 1243.795 ;
    END
  END wd_in[1686]
  PIN wd_in[1687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1243.865 0.070 1243.935 ;
    END
  END wd_in[1687]
  PIN wd_in[1688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1244.005 0.070 1244.075 ;
    END
  END wd_in[1688]
  PIN wd_in[1689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1244.145 0.070 1244.215 ;
    END
  END wd_in[1689]
  PIN wd_in[1690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1244.285 0.070 1244.355 ;
    END
  END wd_in[1690]
  PIN wd_in[1691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1244.425 0.070 1244.495 ;
    END
  END wd_in[1691]
  PIN wd_in[1692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1244.565 0.070 1244.635 ;
    END
  END wd_in[1692]
  PIN wd_in[1693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1244.705 0.070 1244.775 ;
    END
  END wd_in[1693]
  PIN wd_in[1694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1244.845 0.070 1244.915 ;
    END
  END wd_in[1694]
  PIN wd_in[1695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1244.985 0.070 1245.055 ;
    END
  END wd_in[1695]
  PIN wd_in[1696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1245.125 0.070 1245.195 ;
    END
  END wd_in[1696]
  PIN wd_in[1697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1245.265 0.070 1245.335 ;
    END
  END wd_in[1697]
  PIN wd_in[1698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1245.405 0.070 1245.475 ;
    END
  END wd_in[1698]
  PIN wd_in[1699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1245.545 0.070 1245.615 ;
    END
  END wd_in[1699]
  PIN wd_in[1700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1245.685 0.070 1245.755 ;
    END
  END wd_in[1700]
  PIN wd_in[1701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1245.825 0.070 1245.895 ;
    END
  END wd_in[1701]
  PIN wd_in[1702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1245.965 0.070 1246.035 ;
    END
  END wd_in[1702]
  PIN wd_in[1703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1246.105 0.070 1246.175 ;
    END
  END wd_in[1703]
  PIN wd_in[1704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1246.245 0.070 1246.315 ;
    END
  END wd_in[1704]
  PIN wd_in[1705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1246.385 0.070 1246.455 ;
    END
  END wd_in[1705]
  PIN wd_in[1706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1246.525 0.070 1246.595 ;
    END
  END wd_in[1706]
  PIN wd_in[1707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1246.665 0.070 1246.735 ;
    END
  END wd_in[1707]
  PIN wd_in[1708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1246.805 0.070 1246.875 ;
    END
  END wd_in[1708]
  PIN wd_in[1709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1246.945 0.070 1247.015 ;
    END
  END wd_in[1709]
  PIN wd_in[1710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1247.085 0.070 1247.155 ;
    END
  END wd_in[1710]
  PIN wd_in[1711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1247.225 0.070 1247.295 ;
    END
  END wd_in[1711]
  PIN wd_in[1712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1247.365 0.070 1247.435 ;
    END
  END wd_in[1712]
  PIN wd_in[1713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1247.505 0.070 1247.575 ;
    END
  END wd_in[1713]
  PIN wd_in[1714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1247.645 0.070 1247.715 ;
    END
  END wd_in[1714]
  PIN wd_in[1715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1247.785 0.070 1247.855 ;
    END
  END wd_in[1715]
  PIN wd_in[1716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1247.925 0.070 1247.995 ;
    END
  END wd_in[1716]
  PIN wd_in[1717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1248.065 0.070 1248.135 ;
    END
  END wd_in[1717]
  PIN wd_in[1718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1248.205 0.070 1248.275 ;
    END
  END wd_in[1718]
  PIN wd_in[1719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1248.345 0.070 1248.415 ;
    END
  END wd_in[1719]
  PIN wd_in[1720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1248.485 0.070 1248.555 ;
    END
  END wd_in[1720]
  PIN wd_in[1721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1248.625 0.070 1248.695 ;
    END
  END wd_in[1721]
  PIN wd_in[1722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1248.765 0.070 1248.835 ;
    END
  END wd_in[1722]
  PIN wd_in[1723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1248.905 0.070 1248.975 ;
    END
  END wd_in[1723]
  PIN wd_in[1724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1249.045 0.070 1249.115 ;
    END
  END wd_in[1724]
  PIN wd_in[1725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1249.185 0.070 1249.255 ;
    END
  END wd_in[1725]
  PIN wd_in[1726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1249.325 0.070 1249.395 ;
    END
  END wd_in[1726]
  PIN wd_in[1727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1249.465 0.070 1249.535 ;
    END
  END wd_in[1727]
  PIN wd_in[1728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1249.605 0.070 1249.675 ;
    END
  END wd_in[1728]
  PIN wd_in[1729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1249.745 0.070 1249.815 ;
    END
  END wd_in[1729]
  PIN wd_in[1730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1249.885 0.070 1249.955 ;
    END
  END wd_in[1730]
  PIN wd_in[1731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1250.025 0.070 1250.095 ;
    END
  END wd_in[1731]
  PIN wd_in[1732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1250.165 0.070 1250.235 ;
    END
  END wd_in[1732]
  PIN wd_in[1733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1250.305 0.070 1250.375 ;
    END
  END wd_in[1733]
  PIN wd_in[1734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1250.445 0.070 1250.515 ;
    END
  END wd_in[1734]
  PIN wd_in[1735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1250.585 0.070 1250.655 ;
    END
  END wd_in[1735]
  PIN wd_in[1736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1250.725 0.070 1250.795 ;
    END
  END wd_in[1736]
  PIN wd_in[1737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1250.865 0.070 1250.935 ;
    END
  END wd_in[1737]
  PIN wd_in[1738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.005 0.070 1251.075 ;
    END
  END wd_in[1738]
  PIN wd_in[1739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.145 0.070 1251.215 ;
    END
  END wd_in[1739]
  PIN wd_in[1740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.285 0.070 1251.355 ;
    END
  END wd_in[1740]
  PIN wd_in[1741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.425 0.070 1251.495 ;
    END
  END wd_in[1741]
  PIN wd_in[1742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.565 0.070 1251.635 ;
    END
  END wd_in[1742]
  PIN wd_in[1743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.705 0.070 1251.775 ;
    END
  END wd_in[1743]
  PIN wd_in[1744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.845 0.070 1251.915 ;
    END
  END wd_in[1744]
  PIN wd_in[1745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1251.985 0.070 1252.055 ;
    END
  END wd_in[1745]
  PIN wd_in[1746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1252.125 0.070 1252.195 ;
    END
  END wd_in[1746]
  PIN wd_in[1747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1252.265 0.070 1252.335 ;
    END
  END wd_in[1747]
  PIN wd_in[1748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1252.405 0.070 1252.475 ;
    END
  END wd_in[1748]
  PIN wd_in[1749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1252.545 0.070 1252.615 ;
    END
  END wd_in[1749]
  PIN wd_in[1750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1252.685 0.070 1252.755 ;
    END
  END wd_in[1750]
  PIN wd_in[1751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1252.825 0.070 1252.895 ;
    END
  END wd_in[1751]
  PIN wd_in[1752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1252.965 0.070 1253.035 ;
    END
  END wd_in[1752]
  PIN wd_in[1753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1253.105 0.070 1253.175 ;
    END
  END wd_in[1753]
  PIN wd_in[1754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1253.245 0.070 1253.315 ;
    END
  END wd_in[1754]
  PIN wd_in[1755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1253.385 0.070 1253.455 ;
    END
  END wd_in[1755]
  PIN wd_in[1756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1253.525 0.070 1253.595 ;
    END
  END wd_in[1756]
  PIN wd_in[1757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1253.665 0.070 1253.735 ;
    END
  END wd_in[1757]
  PIN wd_in[1758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1253.805 0.070 1253.875 ;
    END
  END wd_in[1758]
  PIN wd_in[1759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1253.945 0.070 1254.015 ;
    END
  END wd_in[1759]
  PIN wd_in[1760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1254.085 0.070 1254.155 ;
    END
  END wd_in[1760]
  PIN wd_in[1761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1254.225 0.070 1254.295 ;
    END
  END wd_in[1761]
  PIN wd_in[1762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1254.365 0.070 1254.435 ;
    END
  END wd_in[1762]
  PIN wd_in[1763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1254.505 0.070 1254.575 ;
    END
  END wd_in[1763]
  PIN wd_in[1764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1254.645 0.070 1254.715 ;
    END
  END wd_in[1764]
  PIN wd_in[1765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1254.785 0.070 1254.855 ;
    END
  END wd_in[1765]
  PIN wd_in[1766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1254.925 0.070 1254.995 ;
    END
  END wd_in[1766]
  PIN wd_in[1767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1255.065 0.070 1255.135 ;
    END
  END wd_in[1767]
  PIN wd_in[1768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1255.205 0.070 1255.275 ;
    END
  END wd_in[1768]
  PIN wd_in[1769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1255.345 0.070 1255.415 ;
    END
  END wd_in[1769]
  PIN wd_in[1770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1255.485 0.070 1255.555 ;
    END
  END wd_in[1770]
  PIN wd_in[1771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1255.625 0.070 1255.695 ;
    END
  END wd_in[1771]
  PIN wd_in[1772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1255.765 0.070 1255.835 ;
    END
  END wd_in[1772]
  PIN wd_in[1773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1255.905 0.070 1255.975 ;
    END
  END wd_in[1773]
  PIN wd_in[1774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1256.045 0.070 1256.115 ;
    END
  END wd_in[1774]
  PIN wd_in[1775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1256.185 0.070 1256.255 ;
    END
  END wd_in[1775]
  PIN wd_in[1776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1256.325 0.070 1256.395 ;
    END
  END wd_in[1776]
  PIN wd_in[1777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1256.465 0.070 1256.535 ;
    END
  END wd_in[1777]
  PIN wd_in[1778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1256.605 0.070 1256.675 ;
    END
  END wd_in[1778]
  PIN wd_in[1779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1256.745 0.070 1256.815 ;
    END
  END wd_in[1779]
  PIN wd_in[1780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1256.885 0.070 1256.955 ;
    END
  END wd_in[1780]
  PIN wd_in[1781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1257.025 0.070 1257.095 ;
    END
  END wd_in[1781]
  PIN wd_in[1782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1257.165 0.070 1257.235 ;
    END
  END wd_in[1782]
  PIN wd_in[1783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1257.305 0.070 1257.375 ;
    END
  END wd_in[1783]
  PIN wd_in[1784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1257.445 0.070 1257.515 ;
    END
  END wd_in[1784]
  PIN wd_in[1785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1257.585 0.070 1257.655 ;
    END
  END wd_in[1785]
  PIN wd_in[1786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1257.725 0.070 1257.795 ;
    END
  END wd_in[1786]
  PIN wd_in[1787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1257.865 0.070 1257.935 ;
    END
  END wd_in[1787]
  PIN wd_in[1788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1258.005 0.070 1258.075 ;
    END
  END wd_in[1788]
  PIN wd_in[1789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1258.145 0.070 1258.215 ;
    END
  END wd_in[1789]
  PIN wd_in[1790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1258.285 0.070 1258.355 ;
    END
  END wd_in[1790]
  PIN wd_in[1791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1258.425 0.070 1258.495 ;
    END
  END wd_in[1791]
  PIN wd_in[1792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1258.565 0.070 1258.635 ;
    END
  END wd_in[1792]
  PIN wd_in[1793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1258.705 0.070 1258.775 ;
    END
  END wd_in[1793]
  PIN wd_in[1794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1258.845 0.070 1258.915 ;
    END
  END wd_in[1794]
  PIN wd_in[1795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1258.985 0.070 1259.055 ;
    END
  END wd_in[1795]
  PIN wd_in[1796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1259.125 0.070 1259.195 ;
    END
  END wd_in[1796]
  PIN wd_in[1797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1259.265 0.070 1259.335 ;
    END
  END wd_in[1797]
  PIN wd_in[1798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1259.405 0.070 1259.475 ;
    END
  END wd_in[1798]
  PIN wd_in[1799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1259.545 0.070 1259.615 ;
    END
  END wd_in[1799]
  PIN wd_in[1800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1259.685 0.070 1259.755 ;
    END
  END wd_in[1800]
  PIN wd_in[1801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1259.825 0.070 1259.895 ;
    END
  END wd_in[1801]
  PIN wd_in[1802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1259.965 0.070 1260.035 ;
    END
  END wd_in[1802]
  PIN wd_in[1803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1260.105 0.070 1260.175 ;
    END
  END wd_in[1803]
  PIN wd_in[1804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1260.245 0.070 1260.315 ;
    END
  END wd_in[1804]
  PIN wd_in[1805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1260.385 0.070 1260.455 ;
    END
  END wd_in[1805]
  PIN wd_in[1806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1260.525 0.070 1260.595 ;
    END
  END wd_in[1806]
  PIN wd_in[1807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1260.665 0.070 1260.735 ;
    END
  END wd_in[1807]
  PIN wd_in[1808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1260.805 0.070 1260.875 ;
    END
  END wd_in[1808]
  PIN wd_in[1809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1260.945 0.070 1261.015 ;
    END
  END wd_in[1809]
  PIN wd_in[1810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1261.085 0.070 1261.155 ;
    END
  END wd_in[1810]
  PIN wd_in[1811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1261.225 0.070 1261.295 ;
    END
  END wd_in[1811]
  PIN wd_in[1812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1261.365 0.070 1261.435 ;
    END
  END wd_in[1812]
  PIN wd_in[1813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1261.505 0.070 1261.575 ;
    END
  END wd_in[1813]
  PIN wd_in[1814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1261.645 0.070 1261.715 ;
    END
  END wd_in[1814]
  PIN wd_in[1815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1261.785 0.070 1261.855 ;
    END
  END wd_in[1815]
  PIN wd_in[1816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1261.925 0.070 1261.995 ;
    END
  END wd_in[1816]
  PIN wd_in[1817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1262.065 0.070 1262.135 ;
    END
  END wd_in[1817]
  PIN wd_in[1818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1262.205 0.070 1262.275 ;
    END
  END wd_in[1818]
  PIN wd_in[1819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1262.345 0.070 1262.415 ;
    END
  END wd_in[1819]
  PIN wd_in[1820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1262.485 0.070 1262.555 ;
    END
  END wd_in[1820]
  PIN wd_in[1821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1262.625 0.070 1262.695 ;
    END
  END wd_in[1821]
  PIN wd_in[1822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1262.765 0.070 1262.835 ;
    END
  END wd_in[1822]
  PIN wd_in[1823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1262.905 0.070 1262.975 ;
    END
  END wd_in[1823]
  PIN wd_in[1824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1263.045 0.070 1263.115 ;
    END
  END wd_in[1824]
  PIN wd_in[1825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1263.185 0.070 1263.255 ;
    END
  END wd_in[1825]
  PIN wd_in[1826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1263.325 0.070 1263.395 ;
    END
  END wd_in[1826]
  PIN wd_in[1827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1263.465 0.070 1263.535 ;
    END
  END wd_in[1827]
  PIN wd_in[1828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1263.605 0.070 1263.675 ;
    END
  END wd_in[1828]
  PIN wd_in[1829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1263.745 0.070 1263.815 ;
    END
  END wd_in[1829]
  PIN wd_in[1830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1263.885 0.070 1263.955 ;
    END
  END wd_in[1830]
  PIN wd_in[1831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1264.025 0.070 1264.095 ;
    END
  END wd_in[1831]
  PIN wd_in[1832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1264.165 0.070 1264.235 ;
    END
  END wd_in[1832]
  PIN wd_in[1833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1264.305 0.070 1264.375 ;
    END
  END wd_in[1833]
  PIN wd_in[1834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1264.445 0.070 1264.515 ;
    END
  END wd_in[1834]
  PIN wd_in[1835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1264.585 0.070 1264.655 ;
    END
  END wd_in[1835]
  PIN wd_in[1836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1264.725 0.070 1264.795 ;
    END
  END wd_in[1836]
  PIN wd_in[1837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1264.865 0.070 1264.935 ;
    END
  END wd_in[1837]
  PIN wd_in[1838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1265.005 0.070 1265.075 ;
    END
  END wd_in[1838]
  PIN wd_in[1839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1265.145 0.070 1265.215 ;
    END
  END wd_in[1839]
  PIN wd_in[1840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1265.285 0.070 1265.355 ;
    END
  END wd_in[1840]
  PIN wd_in[1841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1265.425 0.070 1265.495 ;
    END
  END wd_in[1841]
  PIN wd_in[1842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1265.565 0.070 1265.635 ;
    END
  END wd_in[1842]
  PIN wd_in[1843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1265.705 0.070 1265.775 ;
    END
  END wd_in[1843]
  PIN wd_in[1844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1265.845 0.070 1265.915 ;
    END
  END wd_in[1844]
  PIN wd_in[1845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1265.985 0.070 1266.055 ;
    END
  END wd_in[1845]
  PIN wd_in[1846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1266.125 0.070 1266.195 ;
    END
  END wd_in[1846]
  PIN wd_in[1847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1266.265 0.070 1266.335 ;
    END
  END wd_in[1847]
  PIN wd_in[1848]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1266.405 0.070 1266.475 ;
    END
  END wd_in[1848]
  PIN wd_in[1849]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1266.545 0.070 1266.615 ;
    END
  END wd_in[1849]
  PIN wd_in[1850]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1266.685 0.070 1266.755 ;
    END
  END wd_in[1850]
  PIN wd_in[1851]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1266.825 0.070 1266.895 ;
    END
  END wd_in[1851]
  PIN wd_in[1852]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1266.965 0.070 1267.035 ;
    END
  END wd_in[1852]
  PIN wd_in[1853]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1267.105 0.070 1267.175 ;
    END
  END wd_in[1853]
  PIN wd_in[1854]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1267.245 0.070 1267.315 ;
    END
  END wd_in[1854]
  PIN wd_in[1855]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1267.385 0.070 1267.455 ;
    END
  END wd_in[1855]
  PIN wd_in[1856]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1267.525 0.070 1267.595 ;
    END
  END wd_in[1856]
  PIN wd_in[1857]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1267.665 0.070 1267.735 ;
    END
  END wd_in[1857]
  PIN wd_in[1858]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1267.805 0.070 1267.875 ;
    END
  END wd_in[1858]
  PIN wd_in[1859]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1267.945 0.070 1268.015 ;
    END
  END wd_in[1859]
  PIN wd_in[1860]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1268.085 0.070 1268.155 ;
    END
  END wd_in[1860]
  PIN wd_in[1861]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1268.225 0.070 1268.295 ;
    END
  END wd_in[1861]
  PIN wd_in[1862]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1268.365 0.070 1268.435 ;
    END
  END wd_in[1862]
  PIN wd_in[1863]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1268.505 0.070 1268.575 ;
    END
  END wd_in[1863]
  PIN wd_in[1864]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1268.645 0.070 1268.715 ;
    END
  END wd_in[1864]
  PIN wd_in[1865]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1268.785 0.070 1268.855 ;
    END
  END wd_in[1865]
  PIN wd_in[1866]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1268.925 0.070 1268.995 ;
    END
  END wd_in[1866]
  PIN wd_in[1867]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1269.065 0.070 1269.135 ;
    END
  END wd_in[1867]
  PIN wd_in[1868]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1269.205 0.070 1269.275 ;
    END
  END wd_in[1868]
  PIN wd_in[1869]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1269.345 0.070 1269.415 ;
    END
  END wd_in[1869]
  PIN wd_in[1870]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1269.485 0.070 1269.555 ;
    END
  END wd_in[1870]
  PIN wd_in[1871]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1269.625 0.070 1269.695 ;
    END
  END wd_in[1871]
  PIN wd_in[1872]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1269.765 0.070 1269.835 ;
    END
  END wd_in[1872]
  PIN wd_in[1873]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1269.905 0.070 1269.975 ;
    END
  END wd_in[1873]
  PIN wd_in[1874]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1270.045 0.070 1270.115 ;
    END
  END wd_in[1874]
  PIN wd_in[1875]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1270.185 0.070 1270.255 ;
    END
  END wd_in[1875]
  PIN wd_in[1876]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1270.325 0.070 1270.395 ;
    END
  END wd_in[1876]
  PIN wd_in[1877]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1270.465 0.070 1270.535 ;
    END
  END wd_in[1877]
  PIN wd_in[1878]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1270.605 0.070 1270.675 ;
    END
  END wd_in[1878]
  PIN wd_in[1879]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1270.745 0.070 1270.815 ;
    END
  END wd_in[1879]
  PIN wd_in[1880]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1270.885 0.070 1270.955 ;
    END
  END wd_in[1880]
  PIN wd_in[1881]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1271.025 0.070 1271.095 ;
    END
  END wd_in[1881]
  PIN wd_in[1882]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1271.165 0.070 1271.235 ;
    END
  END wd_in[1882]
  PIN wd_in[1883]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1271.305 0.070 1271.375 ;
    END
  END wd_in[1883]
  PIN wd_in[1884]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1271.445 0.070 1271.515 ;
    END
  END wd_in[1884]
  PIN wd_in[1885]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1271.585 0.070 1271.655 ;
    END
  END wd_in[1885]
  PIN wd_in[1886]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1271.725 0.070 1271.795 ;
    END
  END wd_in[1886]
  PIN wd_in[1887]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1271.865 0.070 1271.935 ;
    END
  END wd_in[1887]
  PIN wd_in[1888]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.005 0.070 1272.075 ;
    END
  END wd_in[1888]
  PIN wd_in[1889]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.145 0.070 1272.215 ;
    END
  END wd_in[1889]
  PIN wd_in[1890]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.285 0.070 1272.355 ;
    END
  END wd_in[1890]
  PIN wd_in[1891]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.425 0.070 1272.495 ;
    END
  END wd_in[1891]
  PIN wd_in[1892]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.565 0.070 1272.635 ;
    END
  END wd_in[1892]
  PIN wd_in[1893]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.705 0.070 1272.775 ;
    END
  END wd_in[1893]
  PIN wd_in[1894]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.845 0.070 1272.915 ;
    END
  END wd_in[1894]
  PIN wd_in[1895]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1272.985 0.070 1273.055 ;
    END
  END wd_in[1895]
  PIN wd_in[1896]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1273.125 0.070 1273.195 ;
    END
  END wd_in[1896]
  PIN wd_in[1897]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1273.265 0.070 1273.335 ;
    END
  END wd_in[1897]
  PIN wd_in[1898]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1273.405 0.070 1273.475 ;
    END
  END wd_in[1898]
  PIN wd_in[1899]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1273.545 0.070 1273.615 ;
    END
  END wd_in[1899]
  PIN wd_in[1900]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1273.685 0.070 1273.755 ;
    END
  END wd_in[1900]
  PIN wd_in[1901]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1273.825 0.070 1273.895 ;
    END
  END wd_in[1901]
  PIN wd_in[1902]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1273.965 0.070 1274.035 ;
    END
  END wd_in[1902]
  PIN wd_in[1903]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.105 0.070 1274.175 ;
    END
  END wd_in[1903]
  PIN wd_in[1904]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.245 0.070 1274.315 ;
    END
  END wd_in[1904]
  PIN wd_in[1905]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.385 0.070 1274.455 ;
    END
  END wd_in[1905]
  PIN wd_in[1906]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.525 0.070 1274.595 ;
    END
  END wd_in[1906]
  PIN wd_in[1907]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.665 0.070 1274.735 ;
    END
  END wd_in[1907]
  PIN wd_in[1908]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.805 0.070 1274.875 ;
    END
  END wd_in[1908]
  PIN wd_in[1909]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1274.945 0.070 1275.015 ;
    END
  END wd_in[1909]
  PIN wd_in[1910]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1275.085 0.070 1275.155 ;
    END
  END wd_in[1910]
  PIN wd_in[1911]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1275.225 0.070 1275.295 ;
    END
  END wd_in[1911]
  PIN wd_in[1912]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1275.365 0.070 1275.435 ;
    END
  END wd_in[1912]
  PIN wd_in[1913]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1275.505 0.070 1275.575 ;
    END
  END wd_in[1913]
  PIN wd_in[1914]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1275.645 0.070 1275.715 ;
    END
  END wd_in[1914]
  PIN wd_in[1915]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1275.785 0.070 1275.855 ;
    END
  END wd_in[1915]
  PIN wd_in[1916]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1275.925 0.070 1275.995 ;
    END
  END wd_in[1916]
  PIN wd_in[1917]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1276.065 0.070 1276.135 ;
    END
  END wd_in[1917]
  PIN wd_in[1918]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1276.205 0.070 1276.275 ;
    END
  END wd_in[1918]
  PIN wd_in[1919]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1276.345 0.070 1276.415 ;
    END
  END wd_in[1919]
  PIN wd_in[1920]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1276.485 0.070 1276.555 ;
    END
  END wd_in[1920]
  PIN wd_in[1921]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1276.625 0.070 1276.695 ;
    END
  END wd_in[1921]
  PIN wd_in[1922]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1276.765 0.070 1276.835 ;
    END
  END wd_in[1922]
  PIN wd_in[1923]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1276.905 0.070 1276.975 ;
    END
  END wd_in[1923]
  PIN wd_in[1924]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1277.045 0.070 1277.115 ;
    END
  END wd_in[1924]
  PIN wd_in[1925]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1277.185 0.070 1277.255 ;
    END
  END wd_in[1925]
  PIN wd_in[1926]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1277.325 0.070 1277.395 ;
    END
  END wd_in[1926]
  PIN wd_in[1927]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1277.465 0.070 1277.535 ;
    END
  END wd_in[1927]
  PIN wd_in[1928]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1277.605 0.070 1277.675 ;
    END
  END wd_in[1928]
  PIN wd_in[1929]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1277.745 0.070 1277.815 ;
    END
  END wd_in[1929]
  PIN wd_in[1930]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1277.885 0.070 1277.955 ;
    END
  END wd_in[1930]
  PIN wd_in[1931]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1278.025 0.070 1278.095 ;
    END
  END wd_in[1931]
  PIN wd_in[1932]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1278.165 0.070 1278.235 ;
    END
  END wd_in[1932]
  PIN wd_in[1933]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1278.305 0.070 1278.375 ;
    END
  END wd_in[1933]
  PIN wd_in[1934]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1278.445 0.070 1278.515 ;
    END
  END wd_in[1934]
  PIN wd_in[1935]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1278.585 0.070 1278.655 ;
    END
  END wd_in[1935]
  PIN wd_in[1936]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1278.725 0.070 1278.795 ;
    END
  END wd_in[1936]
  PIN wd_in[1937]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1278.865 0.070 1278.935 ;
    END
  END wd_in[1937]
  PIN wd_in[1938]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1279.005 0.070 1279.075 ;
    END
  END wd_in[1938]
  PIN wd_in[1939]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1279.145 0.070 1279.215 ;
    END
  END wd_in[1939]
  PIN wd_in[1940]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1279.285 0.070 1279.355 ;
    END
  END wd_in[1940]
  PIN wd_in[1941]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1279.425 0.070 1279.495 ;
    END
  END wd_in[1941]
  PIN wd_in[1942]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1279.565 0.070 1279.635 ;
    END
  END wd_in[1942]
  PIN wd_in[1943]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1279.705 0.070 1279.775 ;
    END
  END wd_in[1943]
  PIN wd_in[1944]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1279.845 0.070 1279.915 ;
    END
  END wd_in[1944]
  PIN wd_in[1945]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1279.985 0.070 1280.055 ;
    END
  END wd_in[1945]
  PIN wd_in[1946]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1280.125 0.070 1280.195 ;
    END
  END wd_in[1946]
  PIN wd_in[1947]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1280.265 0.070 1280.335 ;
    END
  END wd_in[1947]
  PIN wd_in[1948]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1280.405 0.070 1280.475 ;
    END
  END wd_in[1948]
  PIN wd_in[1949]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1280.545 0.070 1280.615 ;
    END
  END wd_in[1949]
  PIN wd_in[1950]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1280.685 0.070 1280.755 ;
    END
  END wd_in[1950]
  PIN wd_in[1951]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1280.825 0.070 1280.895 ;
    END
  END wd_in[1951]
  PIN wd_in[1952]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1280.965 0.070 1281.035 ;
    END
  END wd_in[1952]
  PIN wd_in[1953]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1281.105 0.070 1281.175 ;
    END
  END wd_in[1953]
  PIN wd_in[1954]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1281.245 0.070 1281.315 ;
    END
  END wd_in[1954]
  PIN wd_in[1955]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1281.385 0.070 1281.455 ;
    END
  END wd_in[1955]
  PIN wd_in[1956]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1281.525 0.070 1281.595 ;
    END
  END wd_in[1956]
  PIN wd_in[1957]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1281.665 0.070 1281.735 ;
    END
  END wd_in[1957]
  PIN wd_in[1958]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1281.805 0.070 1281.875 ;
    END
  END wd_in[1958]
  PIN wd_in[1959]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1281.945 0.070 1282.015 ;
    END
  END wd_in[1959]
  PIN wd_in[1960]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1282.085 0.070 1282.155 ;
    END
  END wd_in[1960]
  PIN wd_in[1961]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1282.225 0.070 1282.295 ;
    END
  END wd_in[1961]
  PIN wd_in[1962]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1282.365 0.070 1282.435 ;
    END
  END wd_in[1962]
  PIN wd_in[1963]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1282.505 0.070 1282.575 ;
    END
  END wd_in[1963]
  PIN wd_in[1964]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1282.645 0.070 1282.715 ;
    END
  END wd_in[1964]
  PIN wd_in[1965]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1282.785 0.070 1282.855 ;
    END
  END wd_in[1965]
  PIN wd_in[1966]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1282.925 0.070 1282.995 ;
    END
  END wd_in[1966]
  PIN wd_in[1967]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1283.065 0.070 1283.135 ;
    END
  END wd_in[1967]
  PIN wd_in[1968]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1283.205 0.070 1283.275 ;
    END
  END wd_in[1968]
  PIN wd_in[1969]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1283.345 0.070 1283.415 ;
    END
  END wd_in[1969]
  PIN wd_in[1970]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1283.485 0.070 1283.555 ;
    END
  END wd_in[1970]
  PIN wd_in[1971]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1283.625 0.070 1283.695 ;
    END
  END wd_in[1971]
  PIN wd_in[1972]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1283.765 0.070 1283.835 ;
    END
  END wd_in[1972]
  PIN wd_in[1973]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1283.905 0.070 1283.975 ;
    END
  END wd_in[1973]
  PIN wd_in[1974]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1284.045 0.070 1284.115 ;
    END
  END wd_in[1974]
  PIN wd_in[1975]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1284.185 0.070 1284.255 ;
    END
  END wd_in[1975]
  PIN wd_in[1976]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1284.325 0.070 1284.395 ;
    END
  END wd_in[1976]
  PIN wd_in[1977]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1284.465 0.070 1284.535 ;
    END
  END wd_in[1977]
  PIN wd_in[1978]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1284.605 0.070 1284.675 ;
    END
  END wd_in[1978]
  PIN wd_in[1979]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1284.745 0.070 1284.815 ;
    END
  END wd_in[1979]
  PIN wd_in[1980]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1284.885 0.070 1284.955 ;
    END
  END wd_in[1980]
  PIN wd_in[1981]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1285.025 0.070 1285.095 ;
    END
  END wd_in[1981]
  PIN wd_in[1982]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1285.165 0.070 1285.235 ;
    END
  END wd_in[1982]
  PIN wd_in[1983]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1285.305 0.070 1285.375 ;
    END
  END wd_in[1983]
  PIN wd_in[1984]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1285.445 0.070 1285.515 ;
    END
  END wd_in[1984]
  PIN wd_in[1985]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1285.585 0.070 1285.655 ;
    END
  END wd_in[1985]
  PIN wd_in[1986]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1285.725 0.070 1285.795 ;
    END
  END wd_in[1986]
  PIN wd_in[1987]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1285.865 0.070 1285.935 ;
    END
  END wd_in[1987]
  PIN wd_in[1988]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1286.005 0.070 1286.075 ;
    END
  END wd_in[1988]
  PIN wd_in[1989]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1286.145 0.070 1286.215 ;
    END
  END wd_in[1989]
  PIN wd_in[1990]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1286.285 0.070 1286.355 ;
    END
  END wd_in[1990]
  PIN wd_in[1991]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1286.425 0.070 1286.495 ;
    END
  END wd_in[1991]
  PIN wd_in[1992]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1286.565 0.070 1286.635 ;
    END
  END wd_in[1992]
  PIN wd_in[1993]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1286.705 0.070 1286.775 ;
    END
  END wd_in[1993]
  PIN wd_in[1994]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1286.845 0.070 1286.915 ;
    END
  END wd_in[1994]
  PIN wd_in[1995]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1286.985 0.070 1287.055 ;
    END
  END wd_in[1995]
  PIN wd_in[1996]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1287.125 0.070 1287.195 ;
    END
  END wd_in[1996]
  PIN wd_in[1997]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1287.265 0.070 1287.335 ;
    END
  END wd_in[1997]
  PIN wd_in[1998]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1287.405 0.070 1287.475 ;
    END
  END wd_in[1998]
  PIN wd_in[1999]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1287.545 0.070 1287.615 ;
    END
  END wd_in[1999]
  PIN wd_in[2000]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1287.685 0.070 1287.755 ;
    END
  END wd_in[2000]
  PIN wd_in[2001]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1287.825 0.070 1287.895 ;
    END
  END wd_in[2001]
  PIN wd_in[2002]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1287.965 0.070 1288.035 ;
    END
  END wd_in[2002]
  PIN wd_in[2003]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1288.105 0.070 1288.175 ;
    END
  END wd_in[2003]
  PIN wd_in[2004]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1288.245 0.070 1288.315 ;
    END
  END wd_in[2004]
  PIN wd_in[2005]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1288.385 0.070 1288.455 ;
    END
  END wd_in[2005]
  PIN wd_in[2006]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1288.525 0.070 1288.595 ;
    END
  END wd_in[2006]
  PIN wd_in[2007]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1288.665 0.070 1288.735 ;
    END
  END wd_in[2007]
  PIN wd_in[2008]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1288.805 0.070 1288.875 ;
    END
  END wd_in[2008]
  PIN wd_in[2009]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1288.945 0.070 1289.015 ;
    END
  END wd_in[2009]
  PIN wd_in[2010]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1289.085 0.070 1289.155 ;
    END
  END wd_in[2010]
  PIN wd_in[2011]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1289.225 0.070 1289.295 ;
    END
  END wd_in[2011]
  PIN wd_in[2012]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1289.365 0.070 1289.435 ;
    END
  END wd_in[2012]
  PIN wd_in[2013]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1289.505 0.070 1289.575 ;
    END
  END wd_in[2013]
  PIN wd_in[2014]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1289.645 0.070 1289.715 ;
    END
  END wd_in[2014]
  PIN wd_in[2015]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1289.785 0.070 1289.855 ;
    END
  END wd_in[2015]
  PIN wd_in[2016]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1289.925 0.070 1289.995 ;
    END
  END wd_in[2016]
  PIN wd_in[2017]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1290.065 0.070 1290.135 ;
    END
  END wd_in[2017]
  PIN wd_in[2018]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1290.205 0.070 1290.275 ;
    END
  END wd_in[2018]
  PIN wd_in[2019]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1290.345 0.070 1290.415 ;
    END
  END wd_in[2019]
  PIN wd_in[2020]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1290.485 0.070 1290.555 ;
    END
  END wd_in[2020]
  PIN wd_in[2021]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1290.625 0.070 1290.695 ;
    END
  END wd_in[2021]
  PIN wd_in[2022]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1290.765 0.070 1290.835 ;
    END
  END wd_in[2022]
  PIN wd_in[2023]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1290.905 0.070 1290.975 ;
    END
  END wd_in[2023]
  PIN wd_in[2024]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1291.045 0.070 1291.115 ;
    END
  END wd_in[2024]
  PIN wd_in[2025]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1291.185 0.070 1291.255 ;
    END
  END wd_in[2025]
  PIN wd_in[2026]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1291.325 0.070 1291.395 ;
    END
  END wd_in[2026]
  PIN wd_in[2027]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1291.465 0.070 1291.535 ;
    END
  END wd_in[2027]
  PIN wd_in[2028]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1291.605 0.070 1291.675 ;
    END
  END wd_in[2028]
  PIN wd_in[2029]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1291.745 0.070 1291.815 ;
    END
  END wd_in[2029]
  PIN wd_in[2030]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1291.885 0.070 1291.955 ;
    END
  END wd_in[2030]
  PIN wd_in[2031]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1292.025 0.070 1292.095 ;
    END
  END wd_in[2031]
  PIN wd_in[2032]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1292.165 0.070 1292.235 ;
    END
  END wd_in[2032]
  PIN wd_in[2033]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1292.305 0.070 1292.375 ;
    END
  END wd_in[2033]
  PIN wd_in[2034]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1292.445 0.070 1292.515 ;
    END
  END wd_in[2034]
  PIN wd_in[2035]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1292.585 0.070 1292.655 ;
    END
  END wd_in[2035]
  PIN wd_in[2036]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1292.725 0.070 1292.795 ;
    END
  END wd_in[2036]
  PIN wd_in[2037]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1292.865 0.070 1292.935 ;
    END
  END wd_in[2037]
  PIN wd_in[2038]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1293.005 0.070 1293.075 ;
    END
  END wd_in[2038]
  PIN wd_in[2039]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1293.145 0.070 1293.215 ;
    END
  END wd_in[2039]
  PIN wd_in[2040]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1293.285 0.070 1293.355 ;
    END
  END wd_in[2040]
  PIN wd_in[2041]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1293.425 0.070 1293.495 ;
    END
  END wd_in[2041]
  PIN wd_in[2042]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1293.565 0.070 1293.635 ;
    END
  END wd_in[2042]
  PIN wd_in[2043]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1293.705 0.070 1293.775 ;
    END
  END wd_in[2043]
  PIN wd_in[2044]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1293.845 0.070 1293.915 ;
    END
  END wd_in[2044]
  PIN wd_in[2045]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1293.985 0.070 1294.055 ;
    END
  END wd_in[2045]
  PIN wd_in[2046]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1294.125 0.070 1294.195 ;
    END
  END wd_in[2046]
  PIN wd_in[2047]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1294.265 0.070 1294.335 ;
    END
  END wd_in[2047]
  PIN wd_in[2048]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1294.405 0.070 1294.475 ;
    END
  END wd_in[2048]
  PIN wd_in[2049]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1294.545 0.070 1294.615 ;
    END
  END wd_in[2049]
  PIN wd_in[2050]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1294.685 0.070 1294.755 ;
    END
  END wd_in[2050]
  PIN wd_in[2051]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1294.825 0.070 1294.895 ;
    END
  END wd_in[2051]
  PIN wd_in[2052]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1294.965 0.070 1295.035 ;
    END
  END wd_in[2052]
  PIN wd_in[2053]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1295.105 0.070 1295.175 ;
    END
  END wd_in[2053]
  PIN wd_in[2054]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1295.245 0.070 1295.315 ;
    END
  END wd_in[2054]
  PIN wd_in[2055]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1295.385 0.070 1295.455 ;
    END
  END wd_in[2055]
  PIN wd_in[2056]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1295.525 0.070 1295.595 ;
    END
  END wd_in[2056]
  PIN wd_in[2057]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1295.665 0.070 1295.735 ;
    END
  END wd_in[2057]
  PIN wd_in[2058]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1295.805 0.070 1295.875 ;
    END
  END wd_in[2058]
  PIN wd_in[2059]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1295.945 0.070 1296.015 ;
    END
  END wd_in[2059]
  PIN wd_in[2060]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1296.085 0.070 1296.155 ;
    END
  END wd_in[2060]
  PIN wd_in[2061]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1296.225 0.070 1296.295 ;
    END
  END wd_in[2061]
  PIN wd_in[2062]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1296.365 0.070 1296.435 ;
    END
  END wd_in[2062]
  PIN wd_in[2063]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1296.505 0.070 1296.575 ;
    END
  END wd_in[2063]
  PIN wd_in[2064]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1296.645 0.070 1296.715 ;
    END
  END wd_in[2064]
  PIN wd_in[2065]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1296.785 0.070 1296.855 ;
    END
  END wd_in[2065]
  PIN wd_in[2066]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1296.925 0.070 1296.995 ;
    END
  END wd_in[2066]
  PIN wd_in[2067]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1297.065 0.070 1297.135 ;
    END
  END wd_in[2067]
  PIN wd_in[2068]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1297.205 0.070 1297.275 ;
    END
  END wd_in[2068]
  PIN wd_in[2069]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1297.345 0.070 1297.415 ;
    END
  END wd_in[2069]
  PIN wd_in[2070]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1297.485 0.070 1297.555 ;
    END
  END wd_in[2070]
  PIN wd_in[2071]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1297.625 0.070 1297.695 ;
    END
  END wd_in[2071]
  PIN wd_in[2072]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1297.765 0.070 1297.835 ;
    END
  END wd_in[2072]
  PIN wd_in[2073]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1297.905 0.070 1297.975 ;
    END
  END wd_in[2073]
  PIN wd_in[2074]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1298.045 0.070 1298.115 ;
    END
  END wd_in[2074]
  PIN wd_in[2075]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1298.185 0.070 1298.255 ;
    END
  END wd_in[2075]
  PIN wd_in[2076]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1298.325 0.070 1298.395 ;
    END
  END wd_in[2076]
  PIN wd_in[2077]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1298.465 0.070 1298.535 ;
    END
  END wd_in[2077]
  PIN wd_in[2078]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1298.605 0.070 1298.675 ;
    END
  END wd_in[2078]
  PIN wd_in[2079]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1298.745 0.070 1298.815 ;
    END
  END wd_in[2079]
  PIN wd_in[2080]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1298.885 0.070 1298.955 ;
    END
  END wd_in[2080]
  PIN wd_in[2081]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1299.025 0.070 1299.095 ;
    END
  END wd_in[2081]
  PIN wd_in[2082]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1299.165 0.070 1299.235 ;
    END
  END wd_in[2082]
  PIN wd_in[2083]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1299.305 0.070 1299.375 ;
    END
  END wd_in[2083]
  PIN wd_in[2084]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1299.445 0.070 1299.515 ;
    END
  END wd_in[2084]
  PIN wd_in[2085]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1299.585 0.070 1299.655 ;
    END
  END wd_in[2085]
  PIN wd_in[2086]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1299.725 0.070 1299.795 ;
    END
  END wd_in[2086]
  PIN wd_in[2087]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1299.865 0.070 1299.935 ;
    END
  END wd_in[2087]
  PIN wd_in[2088]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1300.005 0.070 1300.075 ;
    END
  END wd_in[2088]
  PIN wd_in[2089]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1300.145 0.070 1300.215 ;
    END
  END wd_in[2089]
  PIN wd_in[2090]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1300.285 0.070 1300.355 ;
    END
  END wd_in[2090]
  PIN wd_in[2091]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1300.425 0.070 1300.495 ;
    END
  END wd_in[2091]
  PIN wd_in[2092]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1300.565 0.070 1300.635 ;
    END
  END wd_in[2092]
  PIN wd_in[2093]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1300.705 0.070 1300.775 ;
    END
  END wd_in[2093]
  PIN wd_in[2094]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1300.845 0.070 1300.915 ;
    END
  END wd_in[2094]
  PIN wd_in[2095]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1300.985 0.070 1301.055 ;
    END
  END wd_in[2095]
  PIN wd_in[2096]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1301.125 0.070 1301.195 ;
    END
  END wd_in[2096]
  PIN wd_in[2097]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1301.265 0.070 1301.335 ;
    END
  END wd_in[2097]
  PIN wd_in[2098]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1301.405 0.070 1301.475 ;
    END
  END wd_in[2098]
  PIN wd_in[2099]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1301.545 0.070 1301.615 ;
    END
  END wd_in[2099]
  PIN wd_in[2100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1301.685 0.070 1301.755 ;
    END
  END wd_in[2100]
  PIN wd_in[2101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1301.825 0.070 1301.895 ;
    END
  END wd_in[2101]
  PIN wd_in[2102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1301.965 0.070 1302.035 ;
    END
  END wd_in[2102]
  PIN wd_in[2103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1302.105 0.070 1302.175 ;
    END
  END wd_in[2103]
  PIN wd_in[2104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1302.245 0.070 1302.315 ;
    END
  END wd_in[2104]
  PIN wd_in[2105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1302.385 0.070 1302.455 ;
    END
  END wd_in[2105]
  PIN wd_in[2106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1302.525 0.070 1302.595 ;
    END
  END wd_in[2106]
  PIN wd_in[2107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1302.665 0.070 1302.735 ;
    END
  END wd_in[2107]
  PIN wd_in[2108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1302.805 0.070 1302.875 ;
    END
  END wd_in[2108]
  PIN wd_in[2109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1302.945 0.070 1303.015 ;
    END
  END wd_in[2109]
  PIN wd_in[2110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1303.085 0.070 1303.155 ;
    END
  END wd_in[2110]
  PIN wd_in[2111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1303.225 0.070 1303.295 ;
    END
  END wd_in[2111]
  PIN wd_in[2112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1303.365 0.070 1303.435 ;
    END
  END wd_in[2112]
  PIN wd_in[2113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1303.505 0.070 1303.575 ;
    END
  END wd_in[2113]
  PIN wd_in[2114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1303.645 0.070 1303.715 ;
    END
  END wd_in[2114]
  PIN wd_in[2115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1303.785 0.070 1303.855 ;
    END
  END wd_in[2115]
  PIN wd_in[2116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1303.925 0.070 1303.995 ;
    END
  END wd_in[2116]
  PIN wd_in[2117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1304.065 0.070 1304.135 ;
    END
  END wd_in[2117]
  PIN wd_in[2118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1304.205 0.070 1304.275 ;
    END
  END wd_in[2118]
  PIN wd_in[2119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1304.345 0.070 1304.415 ;
    END
  END wd_in[2119]
  PIN wd_in[2120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1304.485 0.070 1304.555 ;
    END
  END wd_in[2120]
  PIN wd_in[2121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1304.625 0.070 1304.695 ;
    END
  END wd_in[2121]
  PIN wd_in[2122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1304.765 0.070 1304.835 ;
    END
  END wd_in[2122]
  PIN wd_in[2123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1304.905 0.070 1304.975 ;
    END
  END wd_in[2123]
  PIN wd_in[2124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1305.045 0.070 1305.115 ;
    END
  END wd_in[2124]
  PIN wd_in[2125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1305.185 0.070 1305.255 ;
    END
  END wd_in[2125]
  PIN wd_in[2126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1305.325 0.070 1305.395 ;
    END
  END wd_in[2126]
  PIN wd_in[2127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1305.465 0.070 1305.535 ;
    END
  END wd_in[2127]
  PIN wd_in[2128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1305.605 0.070 1305.675 ;
    END
  END wd_in[2128]
  PIN wd_in[2129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1305.745 0.070 1305.815 ;
    END
  END wd_in[2129]
  PIN wd_in[2130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1305.885 0.070 1305.955 ;
    END
  END wd_in[2130]
  PIN wd_in[2131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1306.025 0.070 1306.095 ;
    END
  END wd_in[2131]
  PIN wd_in[2132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1306.165 0.070 1306.235 ;
    END
  END wd_in[2132]
  PIN wd_in[2133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1306.305 0.070 1306.375 ;
    END
  END wd_in[2133]
  PIN wd_in[2134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1306.445 0.070 1306.515 ;
    END
  END wd_in[2134]
  PIN wd_in[2135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1306.585 0.070 1306.655 ;
    END
  END wd_in[2135]
  PIN wd_in[2136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1306.725 0.070 1306.795 ;
    END
  END wd_in[2136]
  PIN wd_in[2137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1306.865 0.070 1306.935 ;
    END
  END wd_in[2137]
  PIN wd_in[2138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1307.005 0.070 1307.075 ;
    END
  END wd_in[2138]
  PIN wd_in[2139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1307.145 0.070 1307.215 ;
    END
  END wd_in[2139]
  PIN wd_in[2140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1307.285 0.070 1307.355 ;
    END
  END wd_in[2140]
  PIN wd_in[2141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1307.425 0.070 1307.495 ;
    END
  END wd_in[2141]
  PIN wd_in[2142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1307.565 0.070 1307.635 ;
    END
  END wd_in[2142]
  PIN wd_in[2143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1307.705 0.070 1307.775 ;
    END
  END wd_in[2143]
  PIN wd_in[2144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1307.845 0.070 1307.915 ;
    END
  END wd_in[2144]
  PIN wd_in[2145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1307.985 0.070 1308.055 ;
    END
  END wd_in[2145]
  PIN wd_in[2146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1308.125 0.070 1308.195 ;
    END
  END wd_in[2146]
  PIN wd_in[2147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1308.265 0.070 1308.335 ;
    END
  END wd_in[2147]
  PIN wd_in[2148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1308.405 0.070 1308.475 ;
    END
  END wd_in[2148]
  PIN wd_in[2149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1308.545 0.070 1308.615 ;
    END
  END wd_in[2149]
  PIN wd_in[2150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1308.685 0.070 1308.755 ;
    END
  END wd_in[2150]
  PIN wd_in[2151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1308.825 0.070 1308.895 ;
    END
  END wd_in[2151]
  PIN wd_in[2152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1308.965 0.070 1309.035 ;
    END
  END wd_in[2152]
  PIN wd_in[2153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1309.105 0.070 1309.175 ;
    END
  END wd_in[2153]
  PIN wd_in[2154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1309.245 0.070 1309.315 ;
    END
  END wd_in[2154]
  PIN wd_in[2155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1309.385 0.070 1309.455 ;
    END
  END wd_in[2155]
  PIN wd_in[2156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1309.525 0.070 1309.595 ;
    END
  END wd_in[2156]
  PIN wd_in[2157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1309.665 0.070 1309.735 ;
    END
  END wd_in[2157]
  PIN wd_in[2158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1309.805 0.070 1309.875 ;
    END
  END wd_in[2158]
  PIN wd_in[2159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1309.945 0.070 1310.015 ;
    END
  END wd_in[2159]
  PIN wd_in[2160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1310.085 0.070 1310.155 ;
    END
  END wd_in[2160]
  PIN wd_in[2161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1310.225 0.070 1310.295 ;
    END
  END wd_in[2161]
  PIN wd_in[2162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1310.365 0.070 1310.435 ;
    END
  END wd_in[2162]
  PIN wd_in[2163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1310.505 0.070 1310.575 ;
    END
  END wd_in[2163]
  PIN wd_in[2164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1310.645 0.070 1310.715 ;
    END
  END wd_in[2164]
  PIN wd_in[2165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1310.785 0.070 1310.855 ;
    END
  END wd_in[2165]
  PIN wd_in[2166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1310.925 0.070 1310.995 ;
    END
  END wd_in[2166]
  PIN wd_in[2167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1311.065 0.070 1311.135 ;
    END
  END wd_in[2167]
  PIN wd_in[2168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1311.205 0.070 1311.275 ;
    END
  END wd_in[2168]
  PIN wd_in[2169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1311.345 0.070 1311.415 ;
    END
  END wd_in[2169]
  PIN wd_in[2170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1311.485 0.070 1311.555 ;
    END
  END wd_in[2170]
  PIN wd_in[2171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1311.625 0.070 1311.695 ;
    END
  END wd_in[2171]
  PIN wd_in[2172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1311.765 0.070 1311.835 ;
    END
  END wd_in[2172]
  PIN wd_in[2173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1311.905 0.070 1311.975 ;
    END
  END wd_in[2173]
  PIN wd_in[2174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1312.045 0.070 1312.115 ;
    END
  END wd_in[2174]
  PIN wd_in[2175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1312.185 0.070 1312.255 ;
    END
  END wd_in[2175]
  PIN wd_in[2176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1312.325 0.070 1312.395 ;
    END
  END wd_in[2176]
  PIN wd_in[2177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1312.465 0.070 1312.535 ;
    END
  END wd_in[2177]
  PIN wd_in[2178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1312.605 0.070 1312.675 ;
    END
  END wd_in[2178]
  PIN wd_in[2179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1312.745 0.070 1312.815 ;
    END
  END wd_in[2179]
  PIN wd_in[2180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1312.885 0.070 1312.955 ;
    END
  END wd_in[2180]
  PIN wd_in[2181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1313.025 0.070 1313.095 ;
    END
  END wd_in[2181]
  PIN wd_in[2182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1313.165 0.070 1313.235 ;
    END
  END wd_in[2182]
  PIN wd_in[2183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1313.305 0.070 1313.375 ;
    END
  END wd_in[2183]
  PIN wd_in[2184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1313.445 0.070 1313.515 ;
    END
  END wd_in[2184]
  PIN wd_in[2185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1313.585 0.070 1313.655 ;
    END
  END wd_in[2185]
  PIN wd_in[2186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1313.725 0.070 1313.795 ;
    END
  END wd_in[2186]
  PIN wd_in[2187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1313.865 0.070 1313.935 ;
    END
  END wd_in[2187]
  PIN wd_in[2188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1314.005 0.070 1314.075 ;
    END
  END wd_in[2188]
  PIN wd_in[2189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1314.145 0.070 1314.215 ;
    END
  END wd_in[2189]
  PIN wd_in[2190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1314.285 0.070 1314.355 ;
    END
  END wd_in[2190]
  PIN wd_in[2191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1314.425 0.070 1314.495 ;
    END
  END wd_in[2191]
  PIN wd_in[2192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1314.565 0.070 1314.635 ;
    END
  END wd_in[2192]
  PIN wd_in[2193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1314.705 0.070 1314.775 ;
    END
  END wd_in[2193]
  PIN wd_in[2194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1314.845 0.070 1314.915 ;
    END
  END wd_in[2194]
  PIN wd_in[2195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1314.985 0.070 1315.055 ;
    END
  END wd_in[2195]
  PIN wd_in[2196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1315.125 0.070 1315.195 ;
    END
  END wd_in[2196]
  PIN wd_in[2197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1315.265 0.070 1315.335 ;
    END
  END wd_in[2197]
  PIN wd_in[2198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1315.405 0.070 1315.475 ;
    END
  END wd_in[2198]
  PIN wd_in[2199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1315.545 0.070 1315.615 ;
    END
  END wd_in[2199]
  PIN wd_in[2200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1315.685 0.070 1315.755 ;
    END
  END wd_in[2200]
  PIN wd_in[2201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1315.825 0.070 1315.895 ;
    END
  END wd_in[2201]
  PIN wd_in[2202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1315.965 0.070 1316.035 ;
    END
  END wd_in[2202]
  PIN wd_in[2203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1316.105 0.070 1316.175 ;
    END
  END wd_in[2203]
  PIN wd_in[2204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1316.245 0.070 1316.315 ;
    END
  END wd_in[2204]
  PIN wd_in[2205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1316.385 0.070 1316.455 ;
    END
  END wd_in[2205]
  PIN wd_in[2206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1316.525 0.070 1316.595 ;
    END
  END wd_in[2206]
  PIN wd_in[2207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1316.665 0.070 1316.735 ;
    END
  END wd_in[2207]
  PIN wd_in[2208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1316.805 0.070 1316.875 ;
    END
  END wd_in[2208]
  PIN wd_in[2209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1316.945 0.070 1317.015 ;
    END
  END wd_in[2209]
  PIN wd_in[2210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1317.085 0.070 1317.155 ;
    END
  END wd_in[2210]
  PIN wd_in[2211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1317.225 0.070 1317.295 ;
    END
  END wd_in[2211]
  PIN wd_in[2212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1317.365 0.070 1317.435 ;
    END
  END wd_in[2212]
  PIN wd_in[2213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1317.505 0.070 1317.575 ;
    END
  END wd_in[2213]
  PIN wd_in[2214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1317.645 0.070 1317.715 ;
    END
  END wd_in[2214]
  PIN wd_in[2215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1317.785 0.070 1317.855 ;
    END
  END wd_in[2215]
  PIN wd_in[2216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1317.925 0.070 1317.995 ;
    END
  END wd_in[2216]
  PIN wd_in[2217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1318.065 0.070 1318.135 ;
    END
  END wd_in[2217]
  PIN wd_in[2218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1318.205 0.070 1318.275 ;
    END
  END wd_in[2218]
  PIN wd_in[2219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1318.345 0.070 1318.415 ;
    END
  END wd_in[2219]
  PIN wd_in[2220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1318.485 0.070 1318.555 ;
    END
  END wd_in[2220]
  PIN wd_in[2221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1318.625 0.070 1318.695 ;
    END
  END wd_in[2221]
  PIN wd_in[2222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1318.765 0.070 1318.835 ;
    END
  END wd_in[2222]
  PIN wd_in[2223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1318.905 0.070 1318.975 ;
    END
  END wd_in[2223]
  PIN wd_in[2224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1319.045 0.070 1319.115 ;
    END
  END wd_in[2224]
  PIN wd_in[2225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1319.185 0.070 1319.255 ;
    END
  END wd_in[2225]
  PIN wd_in[2226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1319.325 0.070 1319.395 ;
    END
  END wd_in[2226]
  PIN wd_in[2227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1319.465 0.070 1319.535 ;
    END
  END wd_in[2227]
  PIN wd_in[2228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1319.605 0.070 1319.675 ;
    END
  END wd_in[2228]
  PIN wd_in[2229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1319.745 0.070 1319.815 ;
    END
  END wd_in[2229]
  PIN wd_in[2230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1319.885 0.070 1319.955 ;
    END
  END wd_in[2230]
  PIN wd_in[2231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1320.025 0.070 1320.095 ;
    END
  END wd_in[2231]
  PIN wd_in[2232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1320.165 0.070 1320.235 ;
    END
  END wd_in[2232]
  PIN wd_in[2233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1320.305 0.070 1320.375 ;
    END
  END wd_in[2233]
  PIN wd_in[2234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1320.445 0.070 1320.515 ;
    END
  END wd_in[2234]
  PIN wd_in[2235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1320.585 0.070 1320.655 ;
    END
  END wd_in[2235]
  PIN wd_in[2236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1320.725 0.070 1320.795 ;
    END
  END wd_in[2236]
  PIN wd_in[2237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1320.865 0.070 1320.935 ;
    END
  END wd_in[2237]
  PIN wd_in[2238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1321.005 0.070 1321.075 ;
    END
  END wd_in[2238]
  PIN wd_in[2239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1321.145 0.070 1321.215 ;
    END
  END wd_in[2239]
  PIN wd_in[2240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1321.285 0.070 1321.355 ;
    END
  END wd_in[2240]
  PIN wd_in[2241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1321.425 0.070 1321.495 ;
    END
  END wd_in[2241]
  PIN wd_in[2242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1321.565 0.070 1321.635 ;
    END
  END wd_in[2242]
  PIN wd_in[2243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1321.705 0.070 1321.775 ;
    END
  END wd_in[2243]
  PIN wd_in[2244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1321.845 0.070 1321.915 ;
    END
  END wd_in[2244]
  PIN wd_in[2245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1321.985 0.070 1322.055 ;
    END
  END wd_in[2245]
  PIN wd_in[2246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1322.125 0.070 1322.195 ;
    END
  END wd_in[2246]
  PIN wd_in[2247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1322.265 0.070 1322.335 ;
    END
  END wd_in[2247]
  PIN wd_in[2248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1322.405 0.070 1322.475 ;
    END
  END wd_in[2248]
  PIN wd_in[2249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1322.545 0.070 1322.615 ;
    END
  END wd_in[2249]
  PIN wd_in[2250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1322.685 0.070 1322.755 ;
    END
  END wd_in[2250]
  PIN wd_in[2251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1322.825 0.070 1322.895 ;
    END
  END wd_in[2251]
  PIN wd_in[2252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1322.965 0.070 1323.035 ;
    END
  END wd_in[2252]
  PIN wd_in[2253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1323.105 0.070 1323.175 ;
    END
  END wd_in[2253]
  PIN wd_in[2254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1323.245 0.070 1323.315 ;
    END
  END wd_in[2254]
  PIN wd_in[2255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1323.385 0.070 1323.455 ;
    END
  END wd_in[2255]
  PIN wd_in[2256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1323.525 0.070 1323.595 ;
    END
  END wd_in[2256]
  PIN wd_in[2257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1323.665 0.070 1323.735 ;
    END
  END wd_in[2257]
  PIN wd_in[2258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1323.805 0.070 1323.875 ;
    END
  END wd_in[2258]
  PIN wd_in[2259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1323.945 0.070 1324.015 ;
    END
  END wd_in[2259]
  PIN wd_in[2260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1324.085 0.070 1324.155 ;
    END
  END wd_in[2260]
  PIN wd_in[2261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1324.225 0.070 1324.295 ;
    END
  END wd_in[2261]
  PIN wd_in[2262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1324.365 0.070 1324.435 ;
    END
  END wd_in[2262]
  PIN wd_in[2263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1324.505 0.070 1324.575 ;
    END
  END wd_in[2263]
  PIN wd_in[2264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1324.645 0.070 1324.715 ;
    END
  END wd_in[2264]
  PIN wd_in[2265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1324.785 0.070 1324.855 ;
    END
  END wd_in[2265]
  PIN wd_in[2266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1324.925 0.070 1324.995 ;
    END
  END wd_in[2266]
  PIN wd_in[2267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1325.065 0.070 1325.135 ;
    END
  END wd_in[2267]
  PIN wd_in[2268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1325.205 0.070 1325.275 ;
    END
  END wd_in[2268]
  PIN wd_in[2269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1325.345 0.070 1325.415 ;
    END
  END wd_in[2269]
  PIN wd_in[2270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1325.485 0.070 1325.555 ;
    END
  END wd_in[2270]
  PIN wd_in[2271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1325.625 0.070 1325.695 ;
    END
  END wd_in[2271]
  PIN wd_in[2272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1325.765 0.070 1325.835 ;
    END
  END wd_in[2272]
  PIN wd_in[2273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1325.905 0.070 1325.975 ;
    END
  END wd_in[2273]
  PIN wd_in[2274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1326.045 0.070 1326.115 ;
    END
  END wd_in[2274]
  PIN wd_in[2275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1326.185 0.070 1326.255 ;
    END
  END wd_in[2275]
  PIN wd_in[2276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1326.325 0.070 1326.395 ;
    END
  END wd_in[2276]
  PIN wd_in[2277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1326.465 0.070 1326.535 ;
    END
  END wd_in[2277]
  PIN wd_in[2278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1326.605 0.070 1326.675 ;
    END
  END wd_in[2278]
  PIN wd_in[2279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1326.745 0.070 1326.815 ;
    END
  END wd_in[2279]
  PIN wd_in[2280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1326.885 0.070 1326.955 ;
    END
  END wd_in[2280]
  PIN wd_in[2281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1327.025 0.070 1327.095 ;
    END
  END wd_in[2281]
  PIN wd_in[2282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1327.165 0.070 1327.235 ;
    END
  END wd_in[2282]
  PIN wd_in[2283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1327.305 0.070 1327.375 ;
    END
  END wd_in[2283]
  PIN wd_in[2284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1327.445 0.070 1327.515 ;
    END
  END wd_in[2284]
  PIN wd_in[2285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1327.585 0.070 1327.655 ;
    END
  END wd_in[2285]
  PIN wd_in[2286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1327.725 0.070 1327.795 ;
    END
  END wd_in[2286]
  PIN wd_in[2287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1327.865 0.070 1327.935 ;
    END
  END wd_in[2287]
  PIN wd_in[2288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1328.005 0.070 1328.075 ;
    END
  END wd_in[2288]
  PIN wd_in[2289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1328.145 0.070 1328.215 ;
    END
  END wd_in[2289]
  PIN wd_in[2290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1328.285 0.070 1328.355 ;
    END
  END wd_in[2290]
  PIN wd_in[2291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1328.425 0.070 1328.495 ;
    END
  END wd_in[2291]
  PIN wd_in[2292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1328.565 0.070 1328.635 ;
    END
  END wd_in[2292]
  PIN wd_in[2293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1328.705 0.070 1328.775 ;
    END
  END wd_in[2293]
  PIN wd_in[2294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1328.845 0.070 1328.915 ;
    END
  END wd_in[2294]
  PIN wd_in[2295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1328.985 0.070 1329.055 ;
    END
  END wd_in[2295]
  PIN wd_in[2296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1329.125 0.070 1329.195 ;
    END
  END wd_in[2296]
  PIN wd_in[2297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1329.265 0.070 1329.335 ;
    END
  END wd_in[2297]
  PIN wd_in[2298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1329.405 0.070 1329.475 ;
    END
  END wd_in[2298]
  PIN wd_in[2299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1329.545 0.070 1329.615 ;
    END
  END wd_in[2299]
  PIN wd_in[2300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1329.685 0.070 1329.755 ;
    END
  END wd_in[2300]
  PIN wd_in[2301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1329.825 0.070 1329.895 ;
    END
  END wd_in[2301]
  PIN wd_in[2302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1329.965 0.070 1330.035 ;
    END
  END wd_in[2302]
  PIN wd_in[2303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1330.105 0.070 1330.175 ;
    END
  END wd_in[2303]
  PIN wd_in[2304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1330.245 0.070 1330.315 ;
    END
  END wd_in[2304]
  PIN wd_in[2305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1330.385 0.070 1330.455 ;
    END
  END wd_in[2305]
  PIN wd_in[2306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1330.525 0.070 1330.595 ;
    END
  END wd_in[2306]
  PIN wd_in[2307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1330.665 0.070 1330.735 ;
    END
  END wd_in[2307]
  PIN wd_in[2308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1330.805 0.070 1330.875 ;
    END
  END wd_in[2308]
  PIN wd_in[2309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1330.945 0.070 1331.015 ;
    END
  END wd_in[2309]
  PIN wd_in[2310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1331.085 0.070 1331.155 ;
    END
  END wd_in[2310]
  PIN wd_in[2311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1331.225 0.070 1331.295 ;
    END
  END wd_in[2311]
  PIN wd_in[2312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1331.365 0.070 1331.435 ;
    END
  END wd_in[2312]
  PIN wd_in[2313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1331.505 0.070 1331.575 ;
    END
  END wd_in[2313]
  PIN wd_in[2314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1331.645 0.070 1331.715 ;
    END
  END wd_in[2314]
  PIN wd_in[2315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1331.785 0.070 1331.855 ;
    END
  END wd_in[2315]
  PIN wd_in[2316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1331.925 0.070 1331.995 ;
    END
  END wd_in[2316]
  PIN wd_in[2317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1332.065 0.070 1332.135 ;
    END
  END wd_in[2317]
  PIN wd_in[2318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1332.205 0.070 1332.275 ;
    END
  END wd_in[2318]
  PIN wd_in[2319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1332.345 0.070 1332.415 ;
    END
  END wd_in[2319]
  PIN wd_in[2320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1332.485 0.070 1332.555 ;
    END
  END wd_in[2320]
  PIN wd_in[2321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1332.625 0.070 1332.695 ;
    END
  END wd_in[2321]
  PIN wd_in[2322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1332.765 0.070 1332.835 ;
    END
  END wd_in[2322]
  PIN wd_in[2323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1332.905 0.070 1332.975 ;
    END
  END wd_in[2323]
  PIN wd_in[2324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1333.045 0.070 1333.115 ;
    END
  END wd_in[2324]
  PIN wd_in[2325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1333.185 0.070 1333.255 ;
    END
  END wd_in[2325]
  PIN wd_in[2326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1333.325 0.070 1333.395 ;
    END
  END wd_in[2326]
  PIN wd_in[2327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1333.465 0.070 1333.535 ;
    END
  END wd_in[2327]
  PIN wd_in[2328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1333.605 0.070 1333.675 ;
    END
  END wd_in[2328]
  PIN wd_in[2329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1333.745 0.070 1333.815 ;
    END
  END wd_in[2329]
  PIN wd_in[2330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1333.885 0.070 1333.955 ;
    END
  END wd_in[2330]
  PIN wd_in[2331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1334.025 0.070 1334.095 ;
    END
  END wd_in[2331]
  PIN wd_in[2332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1334.165 0.070 1334.235 ;
    END
  END wd_in[2332]
  PIN wd_in[2333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1334.305 0.070 1334.375 ;
    END
  END wd_in[2333]
  PIN wd_in[2334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1334.445 0.070 1334.515 ;
    END
  END wd_in[2334]
  PIN wd_in[2335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1334.585 0.070 1334.655 ;
    END
  END wd_in[2335]
  PIN wd_in[2336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1334.725 0.070 1334.795 ;
    END
  END wd_in[2336]
  PIN wd_in[2337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1334.865 0.070 1334.935 ;
    END
  END wd_in[2337]
  PIN wd_in[2338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1335.005 0.070 1335.075 ;
    END
  END wd_in[2338]
  PIN wd_in[2339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1335.145 0.070 1335.215 ;
    END
  END wd_in[2339]
  PIN wd_in[2340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1335.285 0.070 1335.355 ;
    END
  END wd_in[2340]
  PIN wd_in[2341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1335.425 0.070 1335.495 ;
    END
  END wd_in[2341]
  PIN wd_in[2342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1335.565 0.070 1335.635 ;
    END
  END wd_in[2342]
  PIN wd_in[2343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1335.705 0.070 1335.775 ;
    END
  END wd_in[2343]
  PIN wd_in[2344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1335.845 0.070 1335.915 ;
    END
  END wd_in[2344]
  PIN wd_in[2345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1335.985 0.070 1336.055 ;
    END
  END wd_in[2345]
  PIN wd_in[2346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1336.125 0.070 1336.195 ;
    END
  END wd_in[2346]
  PIN wd_in[2347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1336.265 0.070 1336.335 ;
    END
  END wd_in[2347]
  PIN wd_in[2348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1336.405 0.070 1336.475 ;
    END
  END wd_in[2348]
  PIN wd_in[2349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1336.545 0.070 1336.615 ;
    END
  END wd_in[2349]
  PIN wd_in[2350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1336.685 0.070 1336.755 ;
    END
  END wd_in[2350]
  PIN wd_in[2351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1336.825 0.070 1336.895 ;
    END
  END wd_in[2351]
  PIN wd_in[2352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1336.965 0.070 1337.035 ;
    END
  END wd_in[2352]
  PIN wd_in[2353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1337.105 0.070 1337.175 ;
    END
  END wd_in[2353]
  PIN wd_in[2354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1337.245 0.070 1337.315 ;
    END
  END wd_in[2354]
  PIN wd_in[2355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1337.385 0.070 1337.455 ;
    END
  END wd_in[2355]
  PIN wd_in[2356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1337.525 0.070 1337.595 ;
    END
  END wd_in[2356]
  PIN wd_in[2357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1337.665 0.070 1337.735 ;
    END
  END wd_in[2357]
  PIN wd_in[2358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1337.805 0.070 1337.875 ;
    END
  END wd_in[2358]
  PIN wd_in[2359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1337.945 0.070 1338.015 ;
    END
  END wd_in[2359]
  PIN wd_in[2360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1338.085 0.070 1338.155 ;
    END
  END wd_in[2360]
  PIN wd_in[2361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1338.225 0.070 1338.295 ;
    END
  END wd_in[2361]
  PIN wd_in[2362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1338.365 0.070 1338.435 ;
    END
  END wd_in[2362]
  PIN wd_in[2363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1338.505 0.070 1338.575 ;
    END
  END wd_in[2363]
  PIN wd_in[2364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1338.645 0.070 1338.715 ;
    END
  END wd_in[2364]
  PIN wd_in[2365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1338.785 0.070 1338.855 ;
    END
  END wd_in[2365]
  PIN wd_in[2366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1338.925 0.070 1338.995 ;
    END
  END wd_in[2366]
  PIN wd_in[2367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1339.065 0.070 1339.135 ;
    END
  END wd_in[2367]
  PIN wd_in[2368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1339.205 0.070 1339.275 ;
    END
  END wd_in[2368]
  PIN wd_in[2369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1339.345 0.070 1339.415 ;
    END
  END wd_in[2369]
  PIN wd_in[2370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1339.485 0.070 1339.555 ;
    END
  END wd_in[2370]
  PIN wd_in[2371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1339.625 0.070 1339.695 ;
    END
  END wd_in[2371]
  PIN wd_in[2372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1339.765 0.070 1339.835 ;
    END
  END wd_in[2372]
  PIN wd_in[2373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1339.905 0.070 1339.975 ;
    END
  END wd_in[2373]
  PIN wd_in[2374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1340.045 0.070 1340.115 ;
    END
  END wd_in[2374]
  PIN wd_in[2375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1340.185 0.070 1340.255 ;
    END
  END wd_in[2375]
  PIN wd_in[2376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1340.325 0.070 1340.395 ;
    END
  END wd_in[2376]
  PIN wd_in[2377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1340.465 0.070 1340.535 ;
    END
  END wd_in[2377]
  PIN wd_in[2378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1340.605 0.070 1340.675 ;
    END
  END wd_in[2378]
  PIN wd_in[2379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1340.745 0.070 1340.815 ;
    END
  END wd_in[2379]
  PIN wd_in[2380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1340.885 0.070 1340.955 ;
    END
  END wd_in[2380]
  PIN wd_in[2381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1341.025 0.070 1341.095 ;
    END
  END wd_in[2381]
  PIN wd_in[2382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1341.165 0.070 1341.235 ;
    END
  END wd_in[2382]
  PIN wd_in[2383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1341.305 0.070 1341.375 ;
    END
  END wd_in[2383]
  PIN wd_in[2384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1341.445 0.070 1341.515 ;
    END
  END wd_in[2384]
  PIN wd_in[2385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1341.585 0.070 1341.655 ;
    END
  END wd_in[2385]
  PIN wd_in[2386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1341.725 0.070 1341.795 ;
    END
  END wd_in[2386]
  PIN wd_in[2387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1341.865 0.070 1341.935 ;
    END
  END wd_in[2387]
  PIN wd_in[2388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1342.005 0.070 1342.075 ;
    END
  END wd_in[2388]
  PIN wd_in[2389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1342.145 0.070 1342.215 ;
    END
  END wd_in[2389]
  PIN wd_in[2390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1342.285 0.070 1342.355 ;
    END
  END wd_in[2390]
  PIN wd_in[2391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1342.425 0.070 1342.495 ;
    END
  END wd_in[2391]
  PIN wd_in[2392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1342.565 0.070 1342.635 ;
    END
  END wd_in[2392]
  PIN wd_in[2393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1342.705 0.070 1342.775 ;
    END
  END wd_in[2393]
  PIN wd_in[2394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1342.845 0.070 1342.915 ;
    END
  END wd_in[2394]
  PIN wd_in[2395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1342.985 0.070 1343.055 ;
    END
  END wd_in[2395]
  PIN wd_in[2396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1343.125 0.070 1343.195 ;
    END
  END wd_in[2396]
  PIN wd_in[2397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1343.265 0.070 1343.335 ;
    END
  END wd_in[2397]
  PIN wd_in[2398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1343.405 0.070 1343.475 ;
    END
  END wd_in[2398]
  PIN wd_in[2399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1343.545 0.070 1343.615 ;
    END
  END wd_in[2399]
  PIN wd_in[2400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1343.685 0.070 1343.755 ;
    END
  END wd_in[2400]
  PIN wd_in[2401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1343.825 0.070 1343.895 ;
    END
  END wd_in[2401]
  PIN wd_in[2402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1343.965 0.070 1344.035 ;
    END
  END wd_in[2402]
  PIN wd_in[2403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1344.105 0.070 1344.175 ;
    END
  END wd_in[2403]
  PIN wd_in[2404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1344.245 0.070 1344.315 ;
    END
  END wd_in[2404]
  PIN wd_in[2405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1344.385 0.070 1344.455 ;
    END
  END wd_in[2405]
  PIN wd_in[2406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1344.525 0.070 1344.595 ;
    END
  END wd_in[2406]
  PIN wd_in[2407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1344.665 0.070 1344.735 ;
    END
  END wd_in[2407]
  PIN wd_in[2408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1344.805 0.070 1344.875 ;
    END
  END wd_in[2408]
  PIN wd_in[2409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1344.945 0.070 1345.015 ;
    END
  END wd_in[2409]
  PIN wd_in[2410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1345.085 0.070 1345.155 ;
    END
  END wd_in[2410]
  PIN wd_in[2411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1345.225 0.070 1345.295 ;
    END
  END wd_in[2411]
  PIN wd_in[2412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1345.365 0.070 1345.435 ;
    END
  END wd_in[2412]
  PIN wd_in[2413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1345.505 0.070 1345.575 ;
    END
  END wd_in[2413]
  PIN wd_in[2414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1345.645 0.070 1345.715 ;
    END
  END wd_in[2414]
  PIN wd_in[2415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1345.785 0.070 1345.855 ;
    END
  END wd_in[2415]
  PIN wd_in[2416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1345.925 0.070 1345.995 ;
    END
  END wd_in[2416]
  PIN wd_in[2417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1346.065 0.070 1346.135 ;
    END
  END wd_in[2417]
  PIN wd_in[2418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1346.205 0.070 1346.275 ;
    END
  END wd_in[2418]
  PIN wd_in[2419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1346.345 0.070 1346.415 ;
    END
  END wd_in[2419]
  PIN wd_in[2420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1346.485 0.070 1346.555 ;
    END
  END wd_in[2420]
  PIN wd_in[2421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1346.625 0.070 1346.695 ;
    END
  END wd_in[2421]
  PIN wd_in[2422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1346.765 0.070 1346.835 ;
    END
  END wd_in[2422]
  PIN wd_in[2423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1346.905 0.070 1346.975 ;
    END
  END wd_in[2423]
  PIN wd_in[2424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1347.045 0.070 1347.115 ;
    END
  END wd_in[2424]
  PIN wd_in[2425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1347.185 0.070 1347.255 ;
    END
  END wd_in[2425]
  PIN wd_in[2426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1347.325 0.070 1347.395 ;
    END
  END wd_in[2426]
  PIN wd_in[2427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1347.465 0.070 1347.535 ;
    END
  END wd_in[2427]
  PIN wd_in[2428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1347.605 0.070 1347.675 ;
    END
  END wd_in[2428]
  PIN wd_in[2429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1347.745 0.070 1347.815 ;
    END
  END wd_in[2429]
  PIN wd_in[2430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1347.885 0.070 1347.955 ;
    END
  END wd_in[2430]
  PIN wd_in[2431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1348.025 0.070 1348.095 ;
    END
  END wd_in[2431]
  PIN wd_in[2432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1348.165 0.070 1348.235 ;
    END
  END wd_in[2432]
  PIN wd_in[2433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1348.305 0.070 1348.375 ;
    END
  END wd_in[2433]
  PIN wd_in[2434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1348.445 0.070 1348.515 ;
    END
  END wd_in[2434]
  PIN wd_in[2435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1348.585 0.070 1348.655 ;
    END
  END wd_in[2435]
  PIN wd_in[2436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1348.725 0.070 1348.795 ;
    END
  END wd_in[2436]
  PIN wd_in[2437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1348.865 0.070 1348.935 ;
    END
  END wd_in[2437]
  PIN wd_in[2438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1349.005 0.070 1349.075 ;
    END
  END wd_in[2438]
  PIN wd_in[2439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1349.145 0.070 1349.215 ;
    END
  END wd_in[2439]
  PIN wd_in[2440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1349.285 0.070 1349.355 ;
    END
  END wd_in[2440]
  PIN wd_in[2441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1349.425 0.070 1349.495 ;
    END
  END wd_in[2441]
  PIN wd_in[2442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1349.565 0.070 1349.635 ;
    END
  END wd_in[2442]
  PIN wd_in[2443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1349.705 0.070 1349.775 ;
    END
  END wd_in[2443]
  PIN wd_in[2444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1349.845 0.070 1349.915 ;
    END
  END wd_in[2444]
  PIN wd_in[2445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1349.985 0.070 1350.055 ;
    END
  END wd_in[2445]
  PIN wd_in[2446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1350.125 0.070 1350.195 ;
    END
  END wd_in[2446]
  PIN wd_in[2447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1350.265 0.070 1350.335 ;
    END
  END wd_in[2447]
  PIN wd_in[2448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1350.405 0.070 1350.475 ;
    END
  END wd_in[2448]
  PIN wd_in[2449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1350.545 0.070 1350.615 ;
    END
  END wd_in[2449]
  PIN wd_in[2450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1350.685 0.070 1350.755 ;
    END
  END wd_in[2450]
  PIN wd_in[2451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1350.825 0.070 1350.895 ;
    END
  END wd_in[2451]
  PIN wd_in[2452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1350.965 0.070 1351.035 ;
    END
  END wd_in[2452]
  PIN wd_in[2453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1351.105 0.070 1351.175 ;
    END
  END wd_in[2453]
  PIN wd_in[2454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1351.245 0.070 1351.315 ;
    END
  END wd_in[2454]
  PIN wd_in[2455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1351.385 0.070 1351.455 ;
    END
  END wd_in[2455]
  PIN wd_in[2456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1351.525 0.070 1351.595 ;
    END
  END wd_in[2456]
  PIN wd_in[2457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1351.665 0.070 1351.735 ;
    END
  END wd_in[2457]
  PIN wd_in[2458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1351.805 0.070 1351.875 ;
    END
  END wd_in[2458]
  PIN wd_in[2459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1351.945 0.070 1352.015 ;
    END
  END wd_in[2459]
  PIN wd_in[2460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1352.085 0.070 1352.155 ;
    END
  END wd_in[2460]
  PIN wd_in[2461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1352.225 0.070 1352.295 ;
    END
  END wd_in[2461]
  PIN wd_in[2462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1352.365 0.070 1352.435 ;
    END
  END wd_in[2462]
  PIN wd_in[2463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1352.505 0.070 1352.575 ;
    END
  END wd_in[2463]
  PIN wd_in[2464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1352.645 0.070 1352.715 ;
    END
  END wd_in[2464]
  PIN wd_in[2465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1352.785 0.070 1352.855 ;
    END
  END wd_in[2465]
  PIN wd_in[2466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1352.925 0.070 1352.995 ;
    END
  END wd_in[2466]
  PIN wd_in[2467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1353.065 0.070 1353.135 ;
    END
  END wd_in[2467]
  PIN wd_in[2468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1353.205 0.070 1353.275 ;
    END
  END wd_in[2468]
  PIN wd_in[2469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1353.345 0.070 1353.415 ;
    END
  END wd_in[2469]
  PIN wd_in[2470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1353.485 0.070 1353.555 ;
    END
  END wd_in[2470]
  PIN wd_in[2471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1353.625 0.070 1353.695 ;
    END
  END wd_in[2471]
  PIN wd_in[2472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1353.765 0.070 1353.835 ;
    END
  END wd_in[2472]
  PIN wd_in[2473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1353.905 0.070 1353.975 ;
    END
  END wd_in[2473]
  PIN wd_in[2474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1354.045 0.070 1354.115 ;
    END
  END wd_in[2474]
  PIN wd_in[2475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1354.185 0.070 1354.255 ;
    END
  END wd_in[2475]
  PIN wd_in[2476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1354.325 0.070 1354.395 ;
    END
  END wd_in[2476]
  PIN wd_in[2477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1354.465 0.070 1354.535 ;
    END
  END wd_in[2477]
  PIN wd_in[2478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1354.605 0.070 1354.675 ;
    END
  END wd_in[2478]
  PIN wd_in[2479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1354.745 0.070 1354.815 ;
    END
  END wd_in[2479]
  PIN wd_in[2480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1354.885 0.070 1354.955 ;
    END
  END wd_in[2480]
  PIN wd_in[2481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1355.025 0.070 1355.095 ;
    END
  END wd_in[2481]
  PIN wd_in[2482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1355.165 0.070 1355.235 ;
    END
  END wd_in[2482]
  PIN wd_in[2483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1355.305 0.070 1355.375 ;
    END
  END wd_in[2483]
  PIN wd_in[2484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1355.445 0.070 1355.515 ;
    END
  END wd_in[2484]
  PIN wd_in[2485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1355.585 0.070 1355.655 ;
    END
  END wd_in[2485]
  PIN wd_in[2486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1355.725 0.070 1355.795 ;
    END
  END wd_in[2486]
  PIN wd_in[2487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1355.865 0.070 1355.935 ;
    END
  END wd_in[2487]
  PIN wd_in[2488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1356.005 0.070 1356.075 ;
    END
  END wd_in[2488]
  PIN wd_in[2489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1356.145 0.070 1356.215 ;
    END
  END wd_in[2489]
  PIN wd_in[2490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1356.285 0.070 1356.355 ;
    END
  END wd_in[2490]
  PIN wd_in[2491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1356.425 0.070 1356.495 ;
    END
  END wd_in[2491]
  PIN wd_in[2492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1356.565 0.070 1356.635 ;
    END
  END wd_in[2492]
  PIN wd_in[2493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1356.705 0.070 1356.775 ;
    END
  END wd_in[2493]
  PIN wd_in[2494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1356.845 0.070 1356.915 ;
    END
  END wd_in[2494]
  PIN wd_in[2495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1356.985 0.070 1357.055 ;
    END
  END wd_in[2495]
  PIN wd_in[2496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1357.125 0.070 1357.195 ;
    END
  END wd_in[2496]
  PIN wd_in[2497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1357.265 0.070 1357.335 ;
    END
  END wd_in[2497]
  PIN wd_in[2498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1357.405 0.070 1357.475 ;
    END
  END wd_in[2498]
  PIN wd_in[2499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1357.545 0.070 1357.615 ;
    END
  END wd_in[2499]
  PIN wd_in[2500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1357.685 0.070 1357.755 ;
    END
  END wd_in[2500]
  PIN wd_in[2501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1357.825 0.070 1357.895 ;
    END
  END wd_in[2501]
  PIN wd_in[2502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1357.965 0.070 1358.035 ;
    END
  END wd_in[2502]
  PIN wd_in[2503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1358.105 0.070 1358.175 ;
    END
  END wd_in[2503]
  PIN wd_in[2504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1358.245 0.070 1358.315 ;
    END
  END wd_in[2504]
  PIN wd_in[2505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1358.385 0.070 1358.455 ;
    END
  END wd_in[2505]
  PIN wd_in[2506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1358.525 0.070 1358.595 ;
    END
  END wd_in[2506]
  PIN wd_in[2507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1358.665 0.070 1358.735 ;
    END
  END wd_in[2507]
  PIN wd_in[2508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1358.805 0.070 1358.875 ;
    END
  END wd_in[2508]
  PIN wd_in[2509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1358.945 0.070 1359.015 ;
    END
  END wd_in[2509]
  PIN wd_in[2510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1359.085 0.070 1359.155 ;
    END
  END wd_in[2510]
  PIN wd_in[2511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1359.225 0.070 1359.295 ;
    END
  END wd_in[2511]
  PIN wd_in[2512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1359.365 0.070 1359.435 ;
    END
  END wd_in[2512]
  PIN wd_in[2513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1359.505 0.070 1359.575 ;
    END
  END wd_in[2513]
  PIN wd_in[2514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1359.645 0.070 1359.715 ;
    END
  END wd_in[2514]
  PIN wd_in[2515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1359.785 0.070 1359.855 ;
    END
  END wd_in[2515]
  PIN wd_in[2516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1359.925 0.070 1359.995 ;
    END
  END wd_in[2516]
  PIN wd_in[2517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1360.065 0.070 1360.135 ;
    END
  END wd_in[2517]
  PIN wd_in[2518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1360.205 0.070 1360.275 ;
    END
  END wd_in[2518]
  PIN wd_in[2519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1360.345 0.070 1360.415 ;
    END
  END wd_in[2519]
  PIN wd_in[2520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1360.485 0.070 1360.555 ;
    END
  END wd_in[2520]
  PIN wd_in[2521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1360.625 0.070 1360.695 ;
    END
  END wd_in[2521]
  PIN wd_in[2522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1360.765 0.070 1360.835 ;
    END
  END wd_in[2522]
  PIN wd_in[2523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1360.905 0.070 1360.975 ;
    END
  END wd_in[2523]
  PIN wd_in[2524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1361.045 0.070 1361.115 ;
    END
  END wd_in[2524]
  PIN wd_in[2525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1361.185 0.070 1361.255 ;
    END
  END wd_in[2525]
  PIN wd_in[2526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1361.325 0.070 1361.395 ;
    END
  END wd_in[2526]
  PIN wd_in[2527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1361.465 0.070 1361.535 ;
    END
  END wd_in[2527]
  PIN wd_in[2528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1361.605 0.070 1361.675 ;
    END
  END wd_in[2528]
  PIN wd_in[2529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1361.745 0.070 1361.815 ;
    END
  END wd_in[2529]
  PIN wd_in[2530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1361.885 0.070 1361.955 ;
    END
  END wd_in[2530]
  PIN wd_in[2531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1362.025 0.070 1362.095 ;
    END
  END wd_in[2531]
  PIN wd_in[2532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1362.165 0.070 1362.235 ;
    END
  END wd_in[2532]
  PIN wd_in[2533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1362.305 0.070 1362.375 ;
    END
  END wd_in[2533]
  PIN wd_in[2534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1362.445 0.070 1362.515 ;
    END
  END wd_in[2534]
  PIN wd_in[2535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1362.585 0.070 1362.655 ;
    END
  END wd_in[2535]
  PIN wd_in[2536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1362.725 0.070 1362.795 ;
    END
  END wd_in[2536]
  PIN wd_in[2537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1362.865 0.070 1362.935 ;
    END
  END wd_in[2537]
  PIN wd_in[2538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1363.005 0.070 1363.075 ;
    END
  END wd_in[2538]
  PIN wd_in[2539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1363.145 0.070 1363.215 ;
    END
  END wd_in[2539]
  PIN wd_in[2540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1363.285 0.070 1363.355 ;
    END
  END wd_in[2540]
  PIN wd_in[2541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1363.425 0.070 1363.495 ;
    END
  END wd_in[2541]
  PIN wd_in[2542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1363.565 0.070 1363.635 ;
    END
  END wd_in[2542]
  PIN wd_in[2543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1363.705 0.070 1363.775 ;
    END
  END wd_in[2543]
  PIN wd_in[2544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1363.845 0.070 1363.915 ;
    END
  END wd_in[2544]
  PIN wd_in[2545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1363.985 0.070 1364.055 ;
    END
  END wd_in[2545]
  PIN wd_in[2546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1364.125 0.070 1364.195 ;
    END
  END wd_in[2546]
  PIN wd_in[2547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1364.265 0.070 1364.335 ;
    END
  END wd_in[2547]
  PIN wd_in[2548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1364.405 0.070 1364.475 ;
    END
  END wd_in[2548]
  PIN wd_in[2549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1364.545 0.070 1364.615 ;
    END
  END wd_in[2549]
  PIN wd_in[2550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1364.685 0.070 1364.755 ;
    END
  END wd_in[2550]
  PIN wd_in[2551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1364.825 0.070 1364.895 ;
    END
  END wd_in[2551]
  PIN wd_in[2552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1364.965 0.070 1365.035 ;
    END
  END wd_in[2552]
  PIN wd_in[2553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1365.105 0.070 1365.175 ;
    END
  END wd_in[2553]
  PIN wd_in[2554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1365.245 0.070 1365.315 ;
    END
  END wd_in[2554]
  PIN wd_in[2555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1365.385 0.070 1365.455 ;
    END
  END wd_in[2555]
  PIN wd_in[2556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1365.525 0.070 1365.595 ;
    END
  END wd_in[2556]
  PIN wd_in[2557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1365.665 0.070 1365.735 ;
    END
  END wd_in[2557]
  PIN wd_in[2558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1365.805 0.070 1365.875 ;
    END
  END wd_in[2558]
  PIN wd_in[2559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1365.945 0.070 1366.015 ;
    END
  END wd_in[2559]
  PIN wd_in[2560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1366.085 0.070 1366.155 ;
    END
  END wd_in[2560]
  PIN wd_in[2561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1366.225 0.070 1366.295 ;
    END
  END wd_in[2561]
  PIN wd_in[2562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1366.365 0.070 1366.435 ;
    END
  END wd_in[2562]
  PIN wd_in[2563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1366.505 0.070 1366.575 ;
    END
  END wd_in[2563]
  PIN wd_in[2564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1366.645 0.070 1366.715 ;
    END
  END wd_in[2564]
  PIN wd_in[2565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1366.785 0.070 1366.855 ;
    END
  END wd_in[2565]
  PIN wd_in[2566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1366.925 0.070 1366.995 ;
    END
  END wd_in[2566]
  PIN wd_in[2567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1367.065 0.070 1367.135 ;
    END
  END wd_in[2567]
  PIN wd_in[2568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1367.205 0.070 1367.275 ;
    END
  END wd_in[2568]
  PIN wd_in[2569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1367.345 0.070 1367.415 ;
    END
  END wd_in[2569]
  PIN wd_in[2570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1367.485 0.070 1367.555 ;
    END
  END wd_in[2570]
  PIN wd_in[2571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1367.625 0.070 1367.695 ;
    END
  END wd_in[2571]
  PIN wd_in[2572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1367.765 0.070 1367.835 ;
    END
  END wd_in[2572]
  PIN wd_in[2573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1367.905 0.070 1367.975 ;
    END
  END wd_in[2573]
  PIN wd_in[2574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1368.045 0.070 1368.115 ;
    END
  END wd_in[2574]
  PIN wd_in[2575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1368.185 0.070 1368.255 ;
    END
  END wd_in[2575]
  PIN wd_in[2576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1368.325 0.070 1368.395 ;
    END
  END wd_in[2576]
  PIN wd_in[2577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1368.465 0.070 1368.535 ;
    END
  END wd_in[2577]
  PIN wd_in[2578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1368.605 0.070 1368.675 ;
    END
  END wd_in[2578]
  PIN wd_in[2579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1368.745 0.070 1368.815 ;
    END
  END wd_in[2579]
  PIN wd_in[2580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1368.885 0.070 1368.955 ;
    END
  END wd_in[2580]
  PIN wd_in[2581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1369.025 0.070 1369.095 ;
    END
  END wd_in[2581]
  PIN wd_in[2582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1369.165 0.070 1369.235 ;
    END
  END wd_in[2582]
  PIN wd_in[2583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1369.305 0.070 1369.375 ;
    END
  END wd_in[2583]
  PIN wd_in[2584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1369.445 0.070 1369.515 ;
    END
  END wd_in[2584]
  PIN wd_in[2585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1369.585 0.070 1369.655 ;
    END
  END wd_in[2585]
  PIN wd_in[2586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1369.725 0.070 1369.795 ;
    END
  END wd_in[2586]
  PIN wd_in[2587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1369.865 0.070 1369.935 ;
    END
  END wd_in[2587]
  PIN wd_in[2588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1370.005 0.070 1370.075 ;
    END
  END wd_in[2588]
  PIN wd_in[2589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1370.145 0.070 1370.215 ;
    END
  END wd_in[2589]
  PIN wd_in[2590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1370.285 0.070 1370.355 ;
    END
  END wd_in[2590]
  PIN wd_in[2591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1370.425 0.070 1370.495 ;
    END
  END wd_in[2591]
  PIN wd_in[2592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1370.565 0.070 1370.635 ;
    END
  END wd_in[2592]
  PIN wd_in[2593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1370.705 0.070 1370.775 ;
    END
  END wd_in[2593]
  PIN wd_in[2594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1370.845 0.070 1370.915 ;
    END
  END wd_in[2594]
  PIN wd_in[2595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1370.985 0.070 1371.055 ;
    END
  END wd_in[2595]
  PIN wd_in[2596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1371.125 0.070 1371.195 ;
    END
  END wd_in[2596]
  PIN wd_in[2597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1371.265 0.070 1371.335 ;
    END
  END wd_in[2597]
  PIN wd_in[2598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1371.405 0.070 1371.475 ;
    END
  END wd_in[2598]
  PIN wd_in[2599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1371.545 0.070 1371.615 ;
    END
  END wd_in[2599]
  PIN wd_in[2600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1371.685 0.070 1371.755 ;
    END
  END wd_in[2600]
  PIN wd_in[2601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1371.825 0.070 1371.895 ;
    END
  END wd_in[2601]
  PIN wd_in[2602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1371.965 0.070 1372.035 ;
    END
  END wd_in[2602]
  PIN wd_in[2603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1372.105 0.070 1372.175 ;
    END
  END wd_in[2603]
  PIN wd_in[2604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1372.245 0.070 1372.315 ;
    END
  END wd_in[2604]
  PIN wd_in[2605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1372.385 0.070 1372.455 ;
    END
  END wd_in[2605]
  PIN wd_in[2606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1372.525 0.070 1372.595 ;
    END
  END wd_in[2606]
  PIN wd_in[2607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1372.665 0.070 1372.735 ;
    END
  END wd_in[2607]
  PIN wd_in[2608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1372.805 0.070 1372.875 ;
    END
  END wd_in[2608]
  PIN wd_in[2609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1372.945 0.070 1373.015 ;
    END
  END wd_in[2609]
  PIN wd_in[2610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1373.085 0.070 1373.155 ;
    END
  END wd_in[2610]
  PIN wd_in[2611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1373.225 0.070 1373.295 ;
    END
  END wd_in[2611]
  PIN wd_in[2612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1373.365 0.070 1373.435 ;
    END
  END wd_in[2612]
  PIN wd_in[2613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1373.505 0.070 1373.575 ;
    END
  END wd_in[2613]
  PIN wd_in[2614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1373.645 0.070 1373.715 ;
    END
  END wd_in[2614]
  PIN wd_in[2615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1373.785 0.070 1373.855 ;
    END
  END wd_in[2615]
  PIN wd_in[2616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1373.925 0.070 1373.995 ;
    END
  END wd_in[2616]
  PIN wd_in[2617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1374.065 0.070 1374.135 ;
    END
  END wd_in[2617]
  PIN wd_in[2618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1374.205 0.070 1374.275 ;
    END
  END wd_in[2618]
  PIN wd_in[2619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1374.345 0.070 1374.415 ;
    END
  END wd_in[2619]
  PIN wd_in[2620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1374.485 0.070 1374.555 ;
    END
  END wd_in[2620]
  PIN wd_in[2621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1374.625 0.070 1374.695 ;
    END
  END wd_in[2621]
  PIN wd_in[2622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1374.765 0.070 1374.835 ;
    END
  END wd_in[2622]
  PIN wd_in[2623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1374.905 0.070 1374.975 ;
    END
  END wd_in[2623]
  PIN wd_in[2624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1375.045 0.070 1375.115 ;
    END
  END wd_in[2624]
  PIN wd_in[2625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1375.185 0.070 1375.255 ;
    END
  END wd_in[2625]
  PIN wd_in[2626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1375.325 0.070 1375.395 ;
    END
  END wd_in[2626]
  PIN wd_in[2627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1375.465 0.070 1375.535 ;
    END
  END wd_in[2627]
  PIN wd_in[2628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1375.605 0.070 1375.675 ;
    END
  END wd_in[2628]
  PIN wd_in[2629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1375.745 0.070 1375.815 ;
    END
  END wd_in[2629]
  PIN wd_in[2630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1375.885 0.070 1375.955 ;
    END
  END wd_in[2630]
  PIN wd_in[2631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1376.025 0.070 1376.095 ;
    END
  END wd_in[2631]
  PIN wd_in[2632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1376.165 0.070 1376.235 ;
    END
  END wd_in[2632]
  PIN wd_in[2633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1376.305 0.070 1376.375 ;
    END
  END wd_in[2633]
  PIN wd_in[2634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1376.445 0.070 1376.515 ;
    END
  END wd_in[2634]
  PIN wd_in[2635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1376.585 0.070 1376.655 ;
    END
  END wd_in[2635]
  PIN wd_in[2636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1376.725 0.070 1376.795 ;
    END
  END wd_in[2636]
  PIN wd_in[2637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1376.865 0.070 1376.935 ;
    END
  END wd_in[2637]
  PIN wd_in[2638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1377.005 0.070 1377.075 ;
    END
  END wd_in[2638]
  PIN wd_in[2639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1377.145 0.070 1377.215 ;
    END
  END wd_in[2639]
  PIN wd_in[2640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1377.285 0.070 1377.355 ;
    END
  END wd_in[2640]
  PIN wd_in[2641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1377.425 0.070 1377.495 ;
    END
  END wd_in[2641]
  PIN wd_in[2642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1377.565 0.070 1377.635 ;
    END
  END wd_in[2642]
  PIN wd_in[2643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1377.705 0.070 1377.775 ;
    END
  END wd_in[2643]
  PIN wd_in[2644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1377.845 0.070 1377.915 ;
    END
  END wd_in[2644]
  PIN wd_in[2645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1377.985 0.070 1378.055 ;
    END
  END wd_in[2645]
  PIN wd_in[2646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1378.125 0.070 1378.195 ;
    END
  END wd_in[2646]
  PIN wd_in[2647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1378.265 0.070 1378.335 ;
    END
  END wd_in[2647]
  PIN wd_in[2648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1378.405 0.070 1378.475 ;
    END
  END wd_in[2648]
  PIN wd_in[2649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1378.545 0.070 1378.615 ;
    END
  END wd_in[2649]
  PIN wd_in[2650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1378.685 0.070 1378.755 ;
    END
  END wd_in[2650]
  PIN wd_in[2651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1378.825 0.070 1378.895 ;
    END
  END wd_in[2651]
  PIN wd_in[2652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1378.965 0.070 1379.035 ;
    END
  END wd_in[2652]
  PIN wd_in[2653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1379.105 0.070 1379.175 ;
    END
  END wd_in[2653]
  PIN wd_in[2654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1379.245 0.070 1379.315 ;
    END
  END wd_in[2654]
  PIN wd_in[2655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1379.385 0.070 1379.455 ;
    END
  END wd_in[2655]
  PIN wd_in[2656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1379.525 0.070 1379.595 ;
    END
  END wd_in[2656]
  PIN wd_in[2657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1379.665 0.070 1379.735 ;
    END
  END wd_in[2657]
  PIN wd_in[2658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1379.805 0.070 1379.875 ;
    END
  END wd_in[2658]
  PIN wd_in[2659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1379.945 0.070 1380.015 ;
    END
  END wd_in[2659]
  PIN wd_in[2660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1380.085 0.070 1380.155 ;
    END
  END wd_in[2660]
  PIN wd_in[2661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1380.225 0.070 1380.295 ;
    END
  END wd_in[2661]
  PIN wd_in[2662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1380.365 0.070 1380.435 ;
    END
  END wd_in[2662]
  PIN wd_in[2663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1380.505 0.070 1380.575 ;
    END
  END wd_in[2663]
  PIN wd_in[2664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1380.645 0.070 1380.715 ;
    END
  END wd_in[2664]
  PIN wd_in[2665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1380.785 0.070 1380.855 ;
    END
  END wd_in[2665]
  PIN wd_in[2666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1380.925 0.070 1380.995 ;
    END
  END wd_in[2666]
  PIN wd_in[2667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1381.065 0.070 1381.135 ;
    END
  END wd_in[2667]
  PIN wd_in[2668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1381.205 0.070 1381.275 ;
    END
  END wd_in[2668]
  PIN wd_in[2669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1381.345 0.070 1381.415 ;
    END
  END wd_in[2669]
  PIN wd_in[2670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1381.485 0.070 1381.555 ;
    END
  END wd_in[2670]
  PIN wd_in[2671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1381.625 0.070 1381.695 ;
    END
  END wd_in[2671]
  PIN wd_in[2672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1381.765 0.070 1381.835 ;
    END
  END wd_in[2672]
  PIN wd_in[2673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1381.905 0.070 1381.975 ;
    END
  END wd_in[2673]
  PIN wd_in[2674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1382.045 0.070 1382.115 ;
    END
  END wd_in[2674]
  PIN wd_in[2675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1382.185 0.070 1382.255 ;
    END
  END wd_in[2675]
  PIN wd_in[2676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1382.325 0.070 1382.395 ;
    END
  END wd_in[2676]
  PIN wd_in[2677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1382.465 0.070 1382.535 ;
    END
  END wd_in[2677]
  PIN wd_in[2678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1382.605 0.070 1382.675 ;
    END
  END wd_in[2678]
  PIN wd_in[2679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1382.745 0.070 1382.815 ;
    END
  END wd_in[2679]
  PIN wd_in[2680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1382.885 0.070 1382.955 ;
    END
  END wd_in[2680]
  PIN wd_in[2681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1383.025 0.070 1383.095 ;
    END
  END wd_in[2681]
  PIN wd_in[2682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1383.165 0.070 1383.235 ;
    END
  END wd_in[2682]
  PIN wd_in[2683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1383.305 0.070 1383.375 ;
    END
  END wd_in[2683]
  PIN wd_in[2684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1383.445 0.070 1383.515 ;
    END
  END wd_in[2684]
  PIN wd_in[2685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1383.585 0.070 1383.655 ;
    END
  END wd_in[2685]
  PIN wd_in[2686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1383.725 0.070 1383.795 ;
    END
  END wd_in[2686]
  PIN wd_in[2687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1383.865 0.070 1383.935 ;
    END
  END wd_in[2687]
  PIN wd_in[2688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1384.005 0.070 1384.075 ;
    END
  END wd_in[2688]
  PIN wd_in[2689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1384.145 0.070 1384.215 ;
    END
  END wd_in[2689]
  PIN wd_in[2690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1384.285 0.070 1384.355 ;
    END
  END wd_in[2690]
  PIN wd_in[2691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1384.425 0.070 1384.495 ;
    END
  END wd_in[2691]
  PIN wd_in[2692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1384.565 0.070 1384.635 ;
    END
  END wd_in[2692]
  PIN wd_in[2693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1384.705 0.070 1384.775 ;
    END
  END wd_in[2693]
  PIN wd_in[2694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1384.845 0.070 1384.915 ;
    END
  END wd_in[2694]
  PIN wd_in[2695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1384.985 0.070 1385.055 ;
    END
  END wd_in[2695]
  PIN wd_in[2696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1385.125 0.070 1385.195 ;
    END
  END wd_in[2696]
  PIN wd_in[2697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1385.265 0.070 1385.335 ;
    END
  END wd_in[2697]
  PIN wd_in[2698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1385.405 0.070 1385.475 ;
    END
  END wd_in[2698]
  PIN wd_in[2699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1385.545 0.070 1385.615 ;
    END
  END wd_in[2699]
  PIN wd_in[2700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1385.685 0.070 1385.755 ;
    END
  END wd_in[2700]
  PIN wd_in[2701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1385.825 0.070 1385.895 ;
    END
  END wd_in[2701]
  PIN wd_in[2702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1385.965 0.070 1386.035 ;
    END
  END wd_in[2702]
  PIN wd_in[2703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1386.105 0.070 1386.175 ;
    END
  END wd_in[2703]
  PIN wd_in[2704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1386.245 0.070 1386.315 ;
    END
  END wd_in[2704]
  PIN wd_in[2705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1386.385 0.070 1386.455 ;
    END
  END wd_in[2705]
  PIN wd_in[2706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1386.525 0.070 1386.595 ;
    END
  END wd_in[2706]
  PIN wd_in[2707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1386.665 0.070 1386.735 ;
    END
  END wd_in[2707]
  PIN wd_in[2708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1386.805 0.070 1386.875 ;
    END
  END wd_in[2708]
  PIN wd_in[2709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1386.945 0.070 1387.015 ;
    END
  END wd_in[2709]
  PIN wd_in[2710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1387.085 0.070 1387.155 ;
    END
  END wd_in[2710]
  PIN wd_in[2711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1387.225 0.070 1387.295 ;
    END
  END wd_in[2711]
  PIN wd_in[2712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1387.365 0.070 1387.435 ;
    END
  END wd_in[2712]
  PIN wd_in[2713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1387.505 0.070 1387.575 ;
    END
  END wd_in[2713]
  PIN wd_in[2714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1387.645 0.070 1387.715 ;
    END
  END wd_in[2714]
  PIN wd_in[2715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1387.785 0.070 1387.855 ;
    END
  END wd_in[2715]
  PIN wd_in[2716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1387.925 0.070 1387.995 ;
    END
  END wd_in[2716]
  PIN wd_in[2717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1388.065 0.070 1388.135 ;
    END
  END wd_in[2717]
  PIN wd_in[2718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1388.205 0.070 1388.275 ;
    END
  END wd_in[2718]
  PIN wd_in[2719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1388.345 0.070 1388.415 ;
    END
  END wd_in[2719]
  PIN wd_in[2720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1388.485 0.070 1388.555 ;
    END
  END wd_in[2720]
  PIN wd_in[2721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1388.625 0.070 1388.695 ;
    END
  END wd_in[2721]
  PIN wd_in[2722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1388.765 0.070 1388.835 ;
    END
  END wd_in[2722]
  PIN wd_in[2723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1388.905 0.070 1388.975 ;
    END
  END wd_in[2723]
  PIN wd_in[2724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1389.045 0.070 1389.115 ;
    END
  END wd_in[2724]
  PIN wd_in[2725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1389.185 0.070 1389.255 ;
    END
  END wd_in[2725]
  PIN wd_in[2726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1389.325 0.070 1389.395 ;
    END
  END wd_in[2726]
  PIN wd_in[2727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1389.465 0.070 1389.535 ;
    END
  END wd_in[2727]
  PIN wd_in[2728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1389.605 0.070 1389.675 ;
    END
  END wd_in[2728]
  PIN wd_in[2729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1389.745 0.070 1389.815 ;
    END
  END wd_in[2729]
  PIN wd_in[2730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1389.885 0.070 1389.955 ;
    END
  END wd_in[2730]
  PIN wd_in[2731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1390.025 0.070 1390.095 ;
    END
  END wd_in[2731]
  PIN wd_in[2732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1390.165 0.070 1390.235 ;
    END
  END wd_in[2732]
  PIN wd_in[2733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1390.305 0.070 1390.375 ;
    END
  END wd_in[2733]
  PIN wd_in[2734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1390.445 0.070 1390.515 ;
    END
  END wd_in[2734]
  PIN wd_in[2735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1390.585 0.070 1390.655 ;
    END
  END wd_in[2735]
  PIN wd_in[2736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1390.725 0.070 1390.795 ;
    END
  END wd_in[2736]
  PIN wd_in[2737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1390.865 0.070 1390.935 ;
    END
  END wd_in[2737]
  PIN wd_in[2738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.005 0.070 1391.075 ;
    END
  END wd_in[2738]
  PIN wd_in[2739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.145 0.070 1391.215 ;
    END
  END wd_in[2739]
  PIN wd_in[2740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.285 0.070 1391.355 ;
    END
  END wd_in[2740]
  PIN wd_in[2741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.425 0.070 1391.495 ;
    END
  END wd_in[2741]
  PIN wd_in[2742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.565 0.070 1391.635 ;
    END
  END wd_in[2742]
  PIN wd_in[2743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.705 0.070 1391.775 ;
    END
  END wd_in[2743]
  PIN wd_in[2744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.845 0.070 1391.915 ;
    END
  END wd_in[2744]
  PIN wd_in[2745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1391.985 0.070 1392.055 ;
    END
  END wd_in[2745]
  PIN wd_in[2746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1392.125 0.070 1392.195 ;
    END
  END wd_in[2746]
  PIN wd_in[2747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1392.265 0.070 1392.335 ;
    END
  END wd_in[2747]
  PIN wd_in[2748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1392.405 0.070 1392.475 ;
    END
  END wd_in[2748]
  PIN wd_in[2749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1392.545 0.070 1392.615 ;
    END
  END wd_in[2749]
  PIN wd_in[2750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1392.685 0.070 1392.755 ;
    END
  END wd_in[2750]
  PIN wd_in[2751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1392.825 0.070 1392.895 ;
    END
  END wd_in[2751]
  PIN wd_in[2752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1392.965 0.070 1393.035 ;
    END
  END wd_in[2752]
  PIN wd_in[2753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1393.105 0.070 1393.175 ;
    END
  END wd_in[2753]
  PIN wd_in[2754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1393.245 0.070 1393.315 ;
    END
  END wd_in[2754]
  PIN wd_in[2755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1393.385 0.070 1393.455 ;
    END
  END wd_in[2755]
  PIN wd_in[2756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1393.525 0.070 1393.595 ;
    END
  END wd_in[2756]
  PIN wd_in[2757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1393.665 0.070 1393.735 ;
    END
  END wd_in[2757]
  PIN wd_in[2758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1393.805 0.070 1393.875 ;
    END
  END wd_in[2758]
  PIN wd_in[2759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1393.945 0.070 1394.015 ;
    END
  END wd_in[2759]
  PIN wd_in[2760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1394.085 0.070 1394.155 ;
    END
  END wd_in[2760]
  PIN wd_in[2761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1394.225 0.070 1394.295 ;
    END
  END wd_in[2761]
  PIN wd_in[2762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1394.365 0.070 1394.435 ;
    END
  END wd_in[2762]
  PIN wd_in[2763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1394.505 0.070 1394.575 ;
    END
  END wd_in[2763]
  PIN wd_in[2764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1394.645 0.070 1394.715 ;
    END
  END wd_in[2764]
  PIN wd_in[2765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1394.785 0.070 1394.855 ;
    END
  END wd_in[2765]
  PIN wd_in[2766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1394.925 0.070 1394.995 ;
    END
  END wd_in[2766]
  PIN wd_in[2767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1395.065 0.070 1395.135 ;
    END
  END wd_in[2767]
  PIN wd_in[2768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1395.205 0.070 1395.275 ;
    END
  END wd_in[2768]
  PIN wd_in[2769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1395.345 0.070 1395.415 ;
    END
  END wd_in[2769]
  PIN wd_in[2770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1395.485 0.070 1395.555 ;
    END
  END wd_in[2770]
  PIN wd_in[2771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1395.625 0.070 1395.695 ;
    END
  END wd_in[2771]
  PIN wd_in[2772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1395.765 0.070 1395.835 ;
    END
  END wd_in[2772]
  PIN wd_in[2773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1395.905 0.070 1395.975 ;
    END
  END wd_in[2773]
  PIN wd_in[2774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1396.045 0.070 1396.115 ;
    END
  END wd_in[2774]
  PIN wd_in[2775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1396.185 0.070 1396.255 ;
    END
  END wd_in[2775]
  PIN wd_in[2776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1396.325 0.070 1396.395 ;
    END
  END wd_in[2776]
  PIN wd_in[2777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1396.465 0.070 1396.535 ;
    END
  END wd_in[2777]
  PIN wd_in[2778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1396.605 0.070 1396.675 ;
    END
  END wd_in[2778]
  PIN wd_in[2779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1396.745 0.070 1396.815 ;
    END
  END wd_in[2779]
  PIN wd_in[2780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1396.885 0.070 1396.955 ;
    END
  END wd_in[2780]
  PIN wd_in[2781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1397.025 0.070 1397.095 ;
    END
  END wd_in[2781]
  PIN wd_in[2782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1397.165 0.070 1397.235 ;
    END
  END wd_in[2782]
  PIN wd_in[2783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1397.305 0.070 1397.375 ;
    END
  END wd_in[2783]
  PIN wd_in[2784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1397.445 0.070 1397.515 ;
    END
  END wd_in[2784]
  PIN wd_in[2785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1397.585 0.070 1397.655 ;
    END
  END wd_in[2785]
  PIN wd_in[2786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1397.725 0.070 1397.795 ;
    END
  END wd_in[2786]
  PIN wd_in[2787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1397.865 0.070 1397.935 ;
    END
  END wd_in[2787]
  PIN wd_in[2788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1398.005 0.070 1398.075 ;
    END
  END wd_in[2788]
  PIN wd_in[2789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1398.145 0.070 1398.215 ;
    END
  END wd_in[2789]
  PIN wd_in[2790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1398.285 0.070 1398.355 ;
    END
  END wd_in[2790]
  PIN wd_in[2791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1398.425 0.070 1398.495 ;
    END
  END wd_in[2791]
  PIN wd_in[2792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1398.565 0.070 1398.635 ;
    END
  END wd_in[2792]
  PIN wd_in[2793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1398.705 0.070 1398.775 ;
    END
  END wd_in[2793]
  PIN wd_in[2794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1398.845 0.070 1398.915 ;
    END
  END wd_in[2794]
  PIN wd_in[2795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1398.985 0.070 1399.055 ;
    END
  END wd_in[2795]
  PIN wd_in[2796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1399.125 0.070 1399.195 ;
    END
  END wd_in[2796]
  PIN wd_in[2797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1399.265 0.070 1399.335 ;
    END
  END wd_in[2797]
  PIN wd_in[2798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1399.405 0.070 1399.475 ;
    END
  END wd_in[2798]
  PIN wd_in[2799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1399.545 0.070 1399.615 ;
    END
  END wd_in[2799]
  PIN wd_in[2800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1399.685 0.070 1399.755 ;
    END
  END wd_in[2800]
  PIN wd_in[2801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1399.825 0.070 1399.895 ;
    END
  END wd_in[2801]
  PIN wd_in[2802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1399.965 0.070 1400.035 ;
    END
  END wd_in[2802]
  PIN wd_in[2803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1400.105 0.070 1400.175 ;
    END
  END wd_in[2803]
  PIN wd_in[2804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1400.245 0.070 1400.315 ;
    END
  END wd_in[2804]
  PIN wd_in[2805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1400.385 0.070 1400.455 ;
    END
  END wd_in[2805]
  PIN wd_in[2806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1400.525 0.070 1400.595 ;
    END
  END wd_in[2806]
  PIN wd_in[2807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1400.665 0.070 1400.735 ;
    END
  END wd_in[2807]
  PIN wd_in[2808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1400.805 0.070 1400.875 ;
    END
  END wd_in[2808]
  PIN wd_in[2809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1400.945 0.070 1401.015 ;
    END
  END wd_in[2809]
  PIN wd_in[2810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1401.085 0.070 1401.155 ;
    END
  END wd_in[2810]
  PIN wd_in[2811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1401.225 0.070 1401.295 ;
    END
  END wd_in[2811]
  PIN wd_in[2812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1401.365 0.070 1401.435 ;
    END
  END wd_in[2812]
  PIN wd_in[2813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1401.505 0.070 1401.575 ;
    END
  END wd_in[2813]
  PIN wd_in[2814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1401.645 0.070 1401.715 ;
    END
  END wd_in[2814]
  PIN wd_in[2815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1401.785 0.070 1401.855 ;
    END
  END wd_in[2815]
  PIN wd_in[2816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1401.925 0.070 1401.995 ;
    END
  END wd_in[2816]
  PIN wd_in[2817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1402.065 0.070 1402.135 ;
    END
  END wd_in[2817]
  PIN wd_in[2818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1402.205 0.070 1402.275 ;
    END
  END wd_in[2818]
  PIN wd_in[2819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1402.345 0.070 1402.415 ;
    END
  END wd_in[2819]
  PIN wd_in[2820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1402.485 0.070 1402.555 ;
    END
  END wd_in[2820]
  PIN wd_in[2821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1402.625 0.070 1402.695 ;
    END
  END wd_in[2821]
  PIN wd_in[2822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1402.765 0.070 1402.835 ;
    END
  END wd_in[2822]
  PIN wd_in[2823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1402.905 0.070 1402.975 ;
    END
  END wd_in[2823]
  PIN wd_in[2824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1403.045 0.070 1403.115 ;
    END
  END wd_in[2824]
  PIN wd_in[2825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1403.185 0.070 1403.255 ;
    END
  END wd_in[2825]
  PIN wd_in[2826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1403.325 0.070 1403.395 ;
    END
  END wd_in[2826]
  PIN wd_in[2827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1403.465 0.070 1403.535 ;
    END
  END wd_in[2827]
  PIN wd_in[2828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1403.605 0.070 1403.675 ;
    END
  END wd_in[2828]
  PIN wd_in[2829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1403.745 0.070 1403.815 ;
    END
  END wd_in[2829]
  PIN wd_in[2830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1403.885 0.070 1403.955 ;
    END
  END wd_in[2830]
  PIN wd_in[2831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1404.025 0.070 1404.095 ;
    END
  END wd_in[2831]
  PIN wd_in[2832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1404.165 0.070 1404.235 ;
    END
  END wd_in[2832]
  PIN wd_in[2833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1404.305 0.070 1404.375 ;
    END
  END wd_in[2833]
  PIN wd_in[2834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1404.445 0.070 1404.515 ;
    END
  END wd_in[2834]
  PIN wd_in[2835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1404.585 0.070 1404.655 ;
    END
  END wd_in[2835]
  PIN wd_in[2836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1404.725 0.070 1404.795 ;
    END
  END wd_in[2836]
  PIN wd_in[2837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1404.865 0.070 1404.935 ;
    END
  END wd_in[2837]
  PIN wd_in[2838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1405.005 0.070 1405.075 ;
    END
  END wd_in[2838]
  PIN wd_in[2839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1405.145 0.070 1405.215 ;
    END
  END wd_in[2839]
  PIN wd_in[2840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1405.285 0.070 1405.355 ;
    END
  END wd_in[2840]
  PIN wd_in[2841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1405.425 0.070 1405.495 ;
    END
  END wd_in[2841]
  PIN wd_in[2842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1405.565 0.070 1405.635 ;
    END
  END wd_in[2842]
  PIN wd_in[2843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1405.705 0.070 1405.775 ;
    END
  END wd_in[2843]
  PIN wd_in[2844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1405.845 0.070 1405.915 ;
    END
  END wd_in[2844]
  PIN wd_in[2845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1405.985 0.070 1406.055 ;
    END
  END wd_in[2845]
  PIN wd_in[2846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1406.125 0.070 1406.195 ;
    END
  END wd_in[2846]
  PIN wd_in[2847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1406.265 0.070 1406.335 ;
    END
  END wd_in[2847]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1510.845 0.070 1510.915 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1510.985 0.070 1511.055 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1511.125 0.070 1511.195 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1511.265 0.070 1511.335 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1511.405 0.070 1511.475 ;
    END
  END addr_in[4]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1615.985 0.070 1616.055 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1616.125 0.070 1616.195 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1616.265 0.070 1616.335 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 1617.000 ;
      RECT 3.500 1.400 3.780 1617.000 ;
      RECT 5.740 1.400 6.020 1617.000 ;
      RECT 7.980 1.400 8.260 1617.000 ;
      RECT 10.220 1.400 10.500 1617.000 ;
      RECT 12.460 1.400 12.740 1617.000 ;
      RECT 14.700 1.400 14.980 1617.000 ;
      RECT 16.940 1.400 17.220 1617.000 ;
      RECT 19.180 1.400 19.460 1617.000 ;
      RECT 21.420 1.400 21.700 1617.000 ;
      RECT 23.660 1.400 23.940 1617.000 ;
      RECT 25.900 1.400 26.180 1617.000 ;
      RECT 28.140 1.400 28.420 1617.000 ;
      RECT 30.380 1.400 30.660 1617.000 ;
      RECT 32.620 1.400 32.900 1617.000 ;
      RECT 34.860 1.400 35.140 1617.000 ;
      RECT 37.100 1.400 37.380 1617.000 ;
      RECT 39.340 1.400 39.620 1617.000 ;
      RECT 41.580 1.400 41.860 1617.000 ;
      RECT 43.820 1.400 44.100 1617.000 ;
      RECT 46.060 1.400 46.340 1617.000 ;
      RECT 48.300 1.400 48.580 1617.000 ;
      RECT 50.540 1.400 50.820 1617.000 ;
      RECT 52.780 1.400 53.060 1617.000 ;
      RECT 55.020 1.400 55.300 1617.000 ;
      RECT 57.260 1.400 57.540 1617.000 ;
      RECT 59.500 1.400 59.780 1617.000 ;
      RECT 61.740 1.400 62.020 1617.000 ;
      RECT 63.980 1.400 64.260 1617.000 ;
      RECT 66.220 1.400 66.500 1617.000 ;
      RECT 68.460 1.400 68.740 1617.000 ;
      RECT 70.700 1.400 70.980 1617.000 ;
      RECT 72.940 1.400 73.220 1617.000 ;
      RECT 75.180 1.400 75.460 1617.000 ;
      RECT 77.420 1.400 77.700 1617.000 ;
      RECT 79.660 1.400 79.940 1617.000 ;
      RECT 81.900 1.400 82.180 1617.000 ;
      RECT 84.140 1.400 84.420 1617.000 ;
      RECT 86.380 1.400 86.660 1617.000 ;
      RECT 88.620 1.400 88.900 1617.000 ;
      RECT 90.860 1.400 91.140 1617.000 ;
      RECT 93.100 1.400 93.380 1617.000 ;
      RECT 95.340 1.400 95.620 1617.000 ;
      RECT 97.580 1.400 97.860 1617.000 ;
      RECT 99.820 1.400 100.100 1617.000 ;
      RECT 102.060 1.400 102.340 1617.000 ;
      RECT 104.300 1.400 104.580 1617.000 ;
      RECT 106.540 1.400 106.820 1617.000 ;
      RECT 108.780 1.400 109.060 1617.000 ;
      RECT 111.020 1.400 111.300 1617.000 ;
      RECT 113.260 1.400 113.540 1617.000 ;
      RECT 115.500 1.400 115.780 1617.000 ;
      RECT 117.740 1.400 118.020 1617.000 ;
      RECT 119.980 1.400 120.260 1617.000 ;
      RECT 122.220 1.400 122.500 1617.000 ;
      RECT 124.460 1.400 124.740 1617.000 ;
      RECT 126.700 1.400 126.980 1617.000 ;
      RECT 128.940 1.400 129.220 1617.000 ;
      RECT 131.180 1.400 131.460 1617.000 ;
      RECT 133.420 1.400 133.700 1617.000 ;
      RECT 135.660 1.400 135.940 1617.000 ;
      RECT 137.900 1.400 138.180 1617.000 ;
      RECT 140.140 1.400 140.420 1617.000 ;
      RECT 142.380 1.400 142.660 1617.000 ;
      RECT 144.620 1.400 144.900 1617.000 ;
      RECT 146.860 1.400 147.140 1617.000 ;
      RECT 149.100 1.400 149.380 1617.000 ;
      RECT 151.340 1.400 151.620 1617.000 ;
      RECT 153.580 1.400 153.860 1617.000 ;
      RECT 155.820 1.400 156.100 1617.000 ;
      RECT 158.060 1.400 158.340 1617.000 ;
      RECT 160.300 1.400 160.580 1617.000 ;
      RECT 162.540 1.400 162.820 1617.000 ;
      RECT 164.780 1.400 165.060 1617.000 ;
      RECT 167.020 1.400 167.300 1617.000 ;
      RECT 169.260 1.400 169.540 1617.000 ;
      RECT 171.500 1.400 171.780 1617.000 ;
      RECT 173.740 1.400 174.020 1617.000 ;
      RECT 175.980 1.400 176.260 1617.000 ;
      RECT 178.220 1.400 178.500 1617.000 ;
      RECT 180.460 1.400 180.740 1617.000 ;
      RECT 182.700 1.400 182.980 1617.000 ;
      RECT 184.940 1.400 185.220 1617.000 ;
      RECT 187.180 1.400 187.460 1617.000 ;
      RECT 189.420 1.400 189.700 1617.000 ;
      RECT 191.660 1.400 191.940 1617.000 ;
      RECT 193.900 1.400 194.180 1617.000 ;
      RECT 196.140 1.400 196.420 1617.000 ;
      RECT 198.380 1.400 198.660 1617.000 ;
      RECT 200.620 1.400 200.900 1617.000 ;
      RECT 202.860 1.400 203.140 1617.000 ;
      RECT 205.100 1.400 205.380 1617.000 ;
      RECT 207.340 1.400 207.620 1617.000 ;
      RECT 209.580 1.400 209.860 1617.000 ;
      RECT 211.820 1.400 212.100 1617.000 ;
      RECT 214.060 1.400 214.340 1617.000 ;
      RECT 216.300 1.400 216.580 1617.000 ;
      RECT 218.540 1.400 218.820 1617.000 ;
      RECT 220.780 1.400 221.060 1617.000 ;
      RECT 223.020 1.400 223.300 1617.000 ;
      RECT 225.260 1.400 225.540 1617.000 ;
      RECT 227.500 1.400 227.780 1617.000 ;
      RECT 229.740 1.400 230.020 1617.000 ;
      RECT 231.980 1.400 232.260 1617.000 ;
      RECT 234.220 1.400 234.500 1617.000 ;
      RECT 236.460 1.400 236.740 1617.000 ;
      RECT 238.700 1.400 238.980 1617.000 ;
      RECT 240.940 1.400 241.220 1617.000 ;
      RECT 243.180 1.400 243.460 1617.000 ;
      RECT 245.420 1.400 245.700 1617.000 ;
      RECT 247.660 1.400 247.940 1617.000 ;
      RECT 249.900 1.400 250.180 1617.000 ;
      RECT 252.140 1.400 252.420 1617.000 ;
      RECT 254.380 1.400 254.660 1617.000 ;
      RECT 256.620 1.400 256.900 1617.000 ;
      RECT 258.860 1.400 259.140 1617.000 ;
      RECT 261.100 1.400 261.380 1617.000 ;
      RECT 263.340 1.400 263.620 1617.000 ;
      RECT 265.580 1.400 265.860 1617.000 ;
      RECT 267.820 1.400 268.100 1617.000 ;
      RECT 270.060 1.400 270.340 1617.000 ;
      RECT 272.300 1.400 272.580 1617.000 ;
      RECT 274.540 1.400 274.820 1617.000 ;
      RECT 276.780 1.400 277.060 1617.000 ;
      RECT 279.020 1.400 279.300 1617.000 ;
      RECT 281.260 1.400 281.540 1617.000 ;
      RECT 283.500 1.400 283.780 1617.000 ;
      RECT 285.740 1.400 286.020 1617.000 ;
      RECT 287.980 1.400 288.260 1617.000 ;
      RECT 290.220 1.400 290.500 1617.000 ;
      RECT 292.460 1.400 292.740 1617.000 ;
      RECT 294.700 1.400 294.980 1617.000 ;
      RECT 296.940 1.400 297.220 1617.000 ;
      RECT 299.180 1.400 299.460 1617.000 ;
      RECT 301.420 1.400 301.700 1617.000 ;
      RECT 303.660 1.400 303.940 1617.000 ;
      RECT 305.900 1.400 306.180 1617.000 ;
      RECT 308.140 1.400 308.420 1617.000 ;
      RECT 310.380 1.400 310.660 1617.000 ;
      RECT 312.620 1.400 312.900 1617.000 ;
      RECT 314.860 1.400 315.140 1617.000 ;
      RECT 317.100 1.400 317.380 1617.000 ;
      RECT 319.340 1.400 319.620 1617.000 ;
      RECT 321.580 1.400 321.860 1617.000 ;
      RECT 323.820 1.400 324.100 1617.000 ;
      RECT 326.060 1.400 326.340 1617.000 ;
      RECT 328.300 1.400 328.580 1617.000 ;
      RECT 330.540 1.400 330.820 1617.000 ;
      RECT 332.780 1.400 333.060 1617.000 ;
      RECT 335.020 1.400 335.300 1617.000 ;
      RECT 337.260 1.400 337.540 1617.000 ;
      RECT 339.500 1.400 339.780 1617.000 ;
      RECT 341.740 1.400 342.020 1617.000 ;
      RECT 343.980 1.400 344.260 1617.000 ;
      RECT 346.220 1.400 346.500 1617.000 ;
      RECT 348.460 1.400 348.740 1617.000 ;
      RECT 350.700 1.400 350.980 1617.000 ;
      RECT 352.940 1.400 353.220 1617.000 ;
      RECT 355.180 1.400 355.460 1617.000 ;
      RECT 357.420 1.400 357.700 1617.000 ;
      RECT 359.660 1.400 359.940 1617.000 ;
      RECT 361.900 1.400 362.180 1617.000 ;
      RECT 364.140 1.400 364.420 1617.000 ;
      RECT 366.380 1.400 366.660 1617.000 ;
      RECT 368.620 1.400 368.900 1617.000 ;
      RECT 370.860 1.400 371.140 1617.000 ;
      RECT 373.100 1.400 373.380 1617.000 ;
      RECT 375.340 1.400 375.620 1617.000 ;
      RECT 377.580 1.400 377.860 1617.000 ;
      RECT 379.820 1.400 380.100 1617.000 ;
      RECT 382.060 1.400 382.340 1617.000 ;
      RECT 384.300 1.400 384.580 1617.000 ;
      RECT 386.540 1.400 386.820 1617.000 ;
      RECT 388.780 1.400 389.060 1617.000 ;
      RECT 391.020 1.400 391.300 1617.000 ;
      RECT 393.260 1.400 393.540 1617.000 ;
      RECT 395.500 1.400 395.780 1617.000 ;
      RECT 397.740 1.400 398.020 1617.000 ;
      RECT 399.980 1.400 400.260 1617.000 ;
      RECT 402.220 1.400 402.500 1617.000 ;
      RECT 404.460 1.400 404.740 1617.000 ;
      RECT 406.700 1.400 406.980 1617.000 ;
      RECT 408.940 1.400 409.220 1617.000 ;
      RECT 411.180 1.400 411.460 1617.000 ;
      RECT 413.420 1.400 413.700 1617.000 ;
      RECT 415.660 1.400 415.940 1617.000 ;
      RECT 417.900 1.400 418.180 1617.000 ;
      RECT 420.140 1.400 420.420 1617.000 ;
      RECT 422.380 1.400 422.660 1617.000 ;
      RECT 424.620 1.400 424.900 1617.000 ;
      RECT 426.860 1.400 427.140 1617.000 ;
      RECT 429.100 1.400 429.380 1617.000 ;
      RECT 431.340 1.400 431.620 1617.000 ;
      RECT 433.580 1.400 433.860 1617.000 ;
      RECT 435.820 1.400 436.100 1617.000 ;
      RECT 438.060 1.400 438.340 1617.000 ;
      RECT 440.300 1.400 440.580 1617.000 ;
      RECT 442.540 1.400 442.820 1617.000 ;
      RECT 444.780 1.400 445.060 1617.000 ;
      RECT 447.020 1.400 447.300 1617.000 ;
      RECT 449.260 1.400 449.540 1617.000 ;
      RECT 451.500 1.400 451.780 1617.000 ;
      RECT 453.740 1.400 454.020 1617.000 ;
      RECT 455.980 1.400 456.260 1617.000 ;
      RECT 458.220 1.400 458.500 1617.000 ;
      RECT 460.460 1.400 460.740 1617.000 ;
      RECT 462.700 1.400 462.980 1617.000 ;
      RECT 464.940 1.400 465.220 1617.000 ;
      RECT 467.180 1.400 467.460 1617.000 ;
      RECT 469.420 1.400 469.700 1617.000 ;
      RECT 471.660 1.400 471.940 1617.000 ;
      RECT 473.900 1.400 474.180 1617.000 ;
      RECT 476.140 1.400 476.420 1617.000 ;
      RECT 478.380 1.400 478.660 1617.000 ;
      RECT 480.620 1.400 480.900 1617.000 ;
      RECT 482.860 1.400 483.140 1617.000 ;
      RECT 485.100 1.400 485.380 1617.000 ;
      RECT 487.340 1.400 487.620 1617.000 ;
      RECT 489.580 1.400 489.860 1617.000 ;
      RECT 491.820 1.400 492.100 1617.000 ;
      RECT 494.060 1.400 494.340 1617.000 ;
      RECT 496.300 1.400 496.580 1617.000 ;
      RECT 498.540 1.400 498.820 1617.000 ;
      RECT 500.780 1.400 501.060 1617.000 ;
      RECT 503.020 1.400 503.300 1617.000 ;
      RECT 505.260 1.400 505.540 1617.000 ;
      RECT 507.500 1.400 507.780 1617.000 ;
      RECT 509.740 1.400 510.020 1617.000 ;
      RECT 511.980 1.400 512.260 1617.000 ;
      RECT 514.220 1.400 514.500 1617.000 ;
      RECT 516.460 1.400 516.740 1617.000 ;
      RECT 518.700 1.400 518.980 1617.000 ;
      RECT 520.940 1.400 521.220 1617.000 ;
      RECT 523.180 1.400 523.460 1617.000 ;
      RECT 525.420 1.400 525.700 1617.000 ;
      RECT 527.660 1.400 527.940 1617.000 ;
      RECT 529.900 1.400 530.180 1617.000 ;
      RECT 532.140 1.400 532.420 1617.000 ;
      RECT 534.380 1.400 534.660 1617.000 ;
      RECT 536.620 1.400 536.900 1617.000 ;
      RECT 538.860 1.400 539.140 1617.000 ;
      RECT 541.100 1.400 541.380 1617.000 ;
      RECT 543.340 1.400 543.620 1617.000 ;
      RECT 545.580 1.400 545.860 1617.000 ;
      RECT 547.820 1.400 548.100 1617.000 ;
      RECT 550.060 1.400 550.340 1617.000 ;
      RECT 552.300 1.400 552.580 1617.000 ;
      RECT 554.540 1.400 554.820 1617.000 ;
      RECT 556.780 1.400 557.060 1617.000 ;
      RECT 559.020 1.400 559.300 1617.000 ;
      RECT 561.260 1.400 561.540 1617.000 ;
      RECT 563.500 1.400 563.780 1617.000 ;
      RECT 565.740 1.400 566.020 1617.000 ;
      RECT 567.980 1.400 568.260 1617.000 ;
      RECT 570.220 1.400 570.500 1617.000 ;
      RECT 572.460 1.400 572.740 1617.000 ;
      RECT 574.700 1.400 574.980 1617.000 ;
      RECT 576.940 1.400 577.220 1617.000 ;
      RECT 579.180 1.400 579.460 1617.000 ;
      RECT 581.420 1.400 581.700 1617.000 ;
      RECT 583.660 1.400 583.940 1617.000 ;
      RECT 585.900 1.400 586.180 1617.000 ;
      RECT 588.140 1.400 588.420 1617.000 ;
      RECT 590.380 1.400 590.660 1617.000 ;
      RECT 592.620 1.400 592.900 1617.000 ;
      RECT 594.860 1.400 595.140 1617.000 ;
      RECT 597.100 1.400 597.380 1617.000 ;
      RECT 599.340 1.400 599.620 1617.000 ;
      RECT 601.580 1.400 601.860 1617.000 ;
      RECT 603.820 1.400 604.100 1617.000 ;
      RECT 606.060 1.400 606.340 1617.000 ;
      RECT 608.300 1.400 608.580 1617.000 ;
      RECT 610.540 1.400 610.820 1617.000 ;
      RECT 612.780 1.400 613.060 1617.000 ;
      RECT 615.020 1.400 615.300 1617.000 ;
      RECT 617.260 1.400 617.540 1617.000 ;
      RECT 619.500 1.400 619.780 1617.000 ;
      RECT 621.740 1.400 622.020 1617.000 ;
      RECT 623.980 1.400 624.260 1617.000 ;
      RECT 626.220 1.400 626.500 1617.000 ;
      RECT 628.460 1.400 628.740 1617.000 ;
      RECT 630.700 1.400 630.980 1617.000 ;
      RECT 632.940 1.400 633.220 1617.000 ;
      RECT 635.180 1.400 635.460 1617.000 ;
      RECT 637.420 1.400 637.700 1617.000 ;
      RECT 639.660 1.400 639.940 1617.000 ;
      RECT 641.900 1.400 642.180 1617.000 ;
      RECT 644.140 1.400 644.420 1617.000 ;
      RECT 646.380 1.400 646.660 1617.000 ;
      RECT 648.620 1.400 648.900 1617.000 ;
      RECT 650.860 1.400 651.140 1617.000 ;
      RECT 653.100 1.400 653.380 1617.000 ;
      RECT 655.340 1.400 655.620 1617.000 ;
      RECT 657.580 1.400 657.860 1617.000 ;
      RECT 659.820 1.400 660.100 1617.000 ;
      RECT 662.060 1.400 662.340 1617.000 ;
      RECT 664.300 1.400 664.580 1617.000 ;
      RECT 666.540 1.400 666.820 1617.000 ;
      RECT 668.780 1.400 669.060 1617.000 ;
      RECT 671.020 1.400 671.300 1617.000 ;
      RECT 673.260 1.400 673.540 1617.000 ;
      RECT 675.500 1.400 675.780 1617.000 ;
      RECT 677.740 1.400 678.020 1617.000 ;
      RECT 679.980 1.400 680.260 1617.000 ;
      RECT 682.220 1.400 682.500 1617.000 ;
      RECT 684.460 1.400 684.740 1617.000 ;
      RECT 686.700 1.400 686.980 1617.000 ;
      RECT 688.940 1.400 689.220 1617.000 ;
      RECT 691.180 1.400 691.460 1617.000 ;
      RECT 693.420 1.400 693.700 1617.000 ;
      RECT 695.660 1.400 695.940 1617.000 ;
      RECT 697.900 1.400 698.180 1617.000 ;
      RECT 700.140 1.400 700.420 1617.000 ;
      RECT 702.380 1.400 702.660 1617.000 ;
      RECT 704.620 1.400 704.900 1617.000 ;
      RECT 706.860 1.400 707.140 1617.000 ;
      RECT 709.100 1.400 709.380 1617.000 ;
      RECT 711.340 1.400 711.620 1617.000 ;
      RECT 713.580 1.400 713.860 1617.000 ;
      RECT 715.820 1.400 716.100 1617.000 ;
      RECT 718.060 1.400 718.340 1617.000 ;
      RECT 720.300 1.400 720.580 1617.000 ;
      RECT 722.540 1.400 722.820 1617.000 ;
      RECT 724.780 1.400 725.060 1617.000 ;
      RECT 727.020 1.400 727.300 1617.000 ;
      RECT 729.260 1.400 729.540 1617.000 ;
      RECT 731.500 1.400 731.780 1617.000 ;
      RECT 733.740 1.400 734.020 1617.000 ;
      RECT 735.980 1.400 736.260 1617.000 ;
      RECT 738.220 1.400 738.500 1617.000 ;
      RECT 740.460 1.400 740.740 1617.000 ;
      RECT 742.700 1.400 742.980 1617.000 ;
      RECT 744.940 1.400 745.220 1617.000 ;
      RECT 747.180 1.400 747.460 1617.000 ;
      RECT 749.420 1.400 749.700 1617.000 ;
      RECT 751.660 1.400 751.940 1617.000 ;
      RECT 753.900 1.400 754.180 1617.000 ;
      RECT 756.140 1.400 756.420 1617.000 ;
      RECT 758.380 1.400 758.660 1617.000 ;
      RECT 760.620 1.400 760.900 1617.000 ;
      RECT 762.860 1.400 763.140 1617.000 ;
      RECT 765.100 1.400 765.380 1617.000 ;
      RECT 767.340 1.400 767.620 1617.000 ;
      RECT 769.580 1.400 769.860 1617.000 ;
      RECT 771.820 1.400 772.100 1617.000 ;
      RECT 774.060 1.400 774.340 1617.000 ;
      RECT 776.300 1.400 776.580 1617.000 ;
      RECT 778.540 1.400 778.820 1617.000 ;
      RECT 780.780 1.400 781.060 1617.000 ;
      RECT 783.020 1.400 783.300 1617.000 ;
      RECT 785.260 1.400 785.540 1617.000 ;
      RECT 787.500 1.400 787.780 1617.000 ;
      RECT 789.740 1.400 790.020 1617.000 ;
      RECT 791.980 1.400 792.260 1617.000 ;
      RECT 794.220 1.400 794.500 1617.000 ;
      RECT 796.460 1.400 796.740 1617.000 ;
      RECT 798.700 1.400 798.980 1617.000 ;
      RECT 800.940 1.400 801.220 1617.000 ;
      RECT 803.180 1.400 803.460 1617.000 ;
      RECT 805.420 1.400 805.700 1617.000 ;
      RECT 807.660 1.400 807.940 1617.000 ;
      RECT 809.900 1.400 810.180 1617.000 ;
      RECT 812.140 1.400 812.420 1617.000 ;
      RECT 814.380 1.400 814.660 1617.000 ;
      RECT 816.620 1.400 816.900 1617.000 ;
      RECT 818.860 1.400 819.140 1617.000 ;
      RECT 821.100 1.400 821.380 1617.000 ;
      RECT 823.340 1.400 823.620 1617.000 ;
      RECT 825.580 1.400 825.860 1617.000 ;
      RECT 827.820 1.400 828.100 1617.000 ;
      RECT 830.060 1.400 830.340 1617.000 ;
      RECT 832.300 1.400 832.580 1617.000 ;
      RECT 834.540 1.400 834.820 1617.000 ;
      RECT 836.780 1.400 837.060 1617.000 ;
      RECT 839.020 1.400 839.300 1617.000 ;
      RECT 841.260 1.400 841.540 1617.000 ;
      RECT 843.500 1.400 843.780 1617.000 ;
      RECT 845.740 1.400 846.020 1617.000 ;
      RECT 847.980 1.400 848.260 1617.000 ;
      RECT 850.220 1.400 850.500 1617.000 ;
      RECT 852.460 1.400 852.740 1617.000 ;
      RECT 854.700 1.400 854.980 1617.000 ;
      RECT 856.940 1.400 857.220 1617.000 ;
      RECT 859.180 1.400 859.460 1617.000 ;
      RECT 861.420 1.400 861.700 1617.000 ;
      RECT 863.660 1.400 863.940 1617.000 ;
      RECT 865.900 1.400 866.180 1617.000 ;
      RECT 868.140 1.400 868.420 1617.000 ;
      RECT 870.380 1.400 870.660 1617.000 ;
      RECT 872.620 1.400 872.900 1617.000 ;
      RECT 874.860 1.400 875.140 1617.000 ;
      RECT 877.100 1.400 877.380 1617.000 ;
      RECT 879.340 1.400 879.620 1617.000 ;
      RECT 881.580 1.400 881.860 1617.000 ;
      RECT 883.820 1.400 884.100 1617.000 ;
      RECT 886.060 1.400 886.340 1617.000 ;
      RECT 888.300 1.400 888.580 1617.000 ;
      RECT 890.540 1.400 890.820 1617.000 ;
      RECT 892.780 1.400 893.060 1617.000 ;
      RECT 895.020 1.400 895.300 1617.000 ;
      RECT 897.260 1.400 897.540 1617.000 ;
      RECT 899.500 1.400 899.780 1617.000 ;
      RECT 901.740 1.400 902.020 1617.000 ;
      RECT 903.980 1.400 904.260 1617.000 ;
      RECT 906.220 1.400 906.500 1617.000 ;
      RECT 908.460 1.400 908.740 1617.000 ;
      RECT 910.700 1.400 910.980 1617.000 ;
      RECT 912.940 1.400 913.220 1617.000 ;
      RECT 915.180 1.400 915.460 1617.000 ;
      RECT 917.420 1.400 917.700 1617.000 ;
      RECT 919.660 1.400 919.940 1617.000 ;
      RECT 921.900 1.400 922.180 1617.000 ;
      RECT 924.140 1.400 924.420 1617.000 ;
      RECT 926.380 1.400 926.660 1617.000 ;
      RECT 928.620 1.400 928.900 1617.000 ;
      RECT 930.860 1.400 931.140 1617.000 ;
      RECT 933.100 1.400 933.380 1617.000 ;
      RECT 935.340 1.400 935.620 1617.000 ;
      RECT 937.580 1.400 937.860 1617.000 ;
      RECT 939.820 1.400 940.100 1617.000 ;
      RECT 942.060 1.400 942.340 1617.000 ;
      RECT 944.300 1.400 944.580 1617.000 ;
      RECT 946.540 1.400 946.820 1617.000 ;
      RECT 948.780 1.400 949.060 1617.000 ;
      RECT 951.020 1.400 951.300 1617.000 ;
      RECT 953.260 1.400 953.540 1617.000 ;
      RECT 955.500 1.400 955.780 1617.000 ;
      RECT 957.740 1.400 958.020 1617.000 ;
      RECT 959.980 1.400 960.260 1617.000 ;
      RECT 962.220 1.400 962.500 1617.000 ;
      RECT 964.460 1.400 964.740 1617.000 ;
      RECT 966.700 1.400 966.980 1617.000 ;
      RECT 968.940 1.400 969.220 1617.000 ;
      RECT 971.180 1.400 971.460 1617.000 ;
      RECT 973.420 1.400 973.700 1617.000 ;
      RECT 975.660 1.400 975.940 1617.000 ;
      RECT 977.900 1.400 978.180 1617.000 ;
      RECT 980.140 1.400 980.420 1617.000 ;
      RECT 982.380 1.400 982.660 1617.000 ;
      RECT 984.620 1.400 984.900 1617.000 ;
      RECT 986.860 1.400 987.140 1617.000 ;
      RECT 989.100 1.400 989.380 1617.000 ;
      RECT 991.340 1.400 991.620 1617.000 ;
      RECT 993.580 1.400 993.860 1617.000 ;
      RECT 995.820 1.400 996.100 1617.000 ;
      RECT 998.060 1.400 998.340 1617.000 ;
      RECT 1000.300 1.400 1000.580 1617.000 ;
      RECT 1002.540 1.400 1002.820 1617.000 ;
      RECT 1004.780 1.400 1005.060 1617.000 ;
      RECT 1007.020 1.400 1007.300 1617.000 ;
      RECT 1009.260 1.400 1009.540 1617.000 ;
      RECT 1011.500 1.400 1011.780 1617.000 ;
      RECT 1013.740 1.400 1014.020 1617.000 ;
      RECT 1015.980 1.400 1016.260 1617.000 ;
      RECT 1018.220 1.400 1018.500 1617.000 ;
      RECT 1020.460 1.400 1020.740 1617.000 ;
      RECT 1022.700 1.400 1022.980 1617.000 ;
      RECT 1024.940 1.400 1025.220 1617.000 ;
      RECT 1027.180 1.400 1027.460 1617.000 ;
      RECT 1029.420 1.400 1029.700 1617.000 ;
      RECT 1031.660 1.400 1031.940 1617.000 ;
      RECT 1033.900 1.400 1034.180 1617.000 ;
      RECT 1036.140 1.400 1036.420 1617.000 ;
      RECT 1038.380 1.400 1038.660 1617.000 ;
      RECT 1040.620 1.400 1040.900 1617.000 ;
      RECT 1042.860 1.400 1043.140 1617.000 ;
      RECT 1045.100 1.400 1045.380 1617.000 ;
      RECT 1047.340 1.400 1047.620 1617.000 ;
      RECT 1049.580 1.400 1049.860 1617.000 ;
      RECT 1051.820 1.400 1052.100 1617.000 ;
      RECT 1054.060 1.400 1054.340 1617.000 ;
      RECT 1056.300 1.400 1056.580 1617.000 ;
      RECT 1058.540 1.400 1058.820 1617.000 ;
      RECT 1060.780 1.400 1061.060 1617.000 ;
      RECT 1063.020 1.400 1063.300 1617.000 ;
      RECT 1065.260 1.400 1065.540 1617.000 ;
      RECT 1067.500 1.400 1067.780 1617.000 ;
      RECT 1069.740 1.400 1070.020 1617.000 ;
      RECT 1071.980 1.400 1072.260 1617.000 ;
      RECT 1074.220 1.400 1074.500 1617.000 ;
      RECT 1076.460 1.400 1076.740 1617.000 ;
      RECT 1078.700 1.400 1078.980 1617.000 ;
      RECT 1080.940 1.400 1081.220 1617.000 ;
      RECT 1083.180 1.400 1083.460 1617.000 ;
      RECT 1085.420 1.400 1085.700 1617.000 ;
      RECT 1087.660 1.400 1087.940 1617.000 ;
      RECT 1089.900 1.400 1090.180 1617.000 ;
      RECT 1092.140 1.400 1092.420 1617.000 ;
      RECT 1094.380 1.400 1094.660 1617.000 ;
      RECT 1096.620 1.400 1096.900 1617.000 ;
      RECT 1098.860 1.400 1099.140 1617.000 ;
      RECT 1101.100 1.400 1101.380 1617.000 ;
      RECT 1103.340 1.400 1103.620 1617.000 ;
      RECT 1105.580 1.400 1105.860 1617.000 ;
      RECT 1107.820 1.400 1108.100 1617.000 ;
      RECT 1110.060 1.400 1110.340 1617.000 ;
      RECT 1112.300 1.400 1112.580 1617.000 ;
      RECT 1114.540 1.400 1114.820 1617.000 ;
      RECT 1116.780 1.400 1117.060 1617.000 ;
      RECT 1119.020 1.400 1119.300 1617.000 ;
      RECT 1121.260 1.400 1121.540 1617.000 ;
      RECT 1123.500 1.400 1123.780 1617.000 ;
      RECT 1125.740 1.400 1126.020 1617.000 ;
      RECT 1127.980 1.400 1128.260 1617.000 ;
      RECT 1130.220 1.400 1130.500 1617.000 ;
      RECT 1132.460 1.400 1132.740 1617.000 ;
      RECT 1134.700 1.400 1134.980 1617.000 ;
      RECT 1136.940 1.400 1137.220 1617.000 ;
      RECT 1139.180 1.400 1139.460 1617.000 ;
      RECT 1141.420 1.400 1141.700 1617.000 ;
      RECT 1143.660 1.400 1143.940 1617.000 ;
      RECT 1145.900 1.400 1146.180 1617.000 ;
      RECT 1148.140 1.400 1148.420 1617.000 ;
      RECT 1150.380 1.400 1150.660 1617.000 ;
      RECT 1152.620 1.400 1152.900 1617.000 ;
      RECT 1154.860 1.400 1155.140 1617.000 ;
      RECT 1157.100 1.400 1157.380 1617.000 ;
      RECT 1159.340 1.400 1159.620 1617.000 ;
      RECT 1161.580 1.400 1161.860 1617.000 ;
      RECT 1163.820 1.400 1164.100 1617.000 ;
      RECT 1166.060 1.400 1166.340 1617.000 ;
      RECT 1168.300 1.400 1168.580 1617.000 ;
      RECT 1170.540 1.400 1170.820 1617.000 ;
      RECT 1172.780 1.400 1173.060 1617.000 ;
      RECT 1175.020 1.400 1175.300 1617.000 ;
      RECT 1177.260 1.400 1177.540 1617.000 ;
      RECT 1179.500 1.400 1179.780 1617.000 ;
      RECT 1181.740 1.400 1182.020 1617.000 ;
      RECT 1183.980 1.400 1184.260 1617.000 ;
      RECT 1186.220 1.400 1186.500 1617.000 ;
      RECT 1188.460 1.400 1188.740 1617.000 ;
      RECT 1190.700 1.400 1190.980 1617.000 ;
      RECT 1192.940 1.400 1193.220 1617.000 ;
      RECT 1195.180 1.400 1195.460 1617.000 ;
      RECT 1197.420 1.400 1197.700 1617.000 ;
      RECT 1199.660 1.400 1199.940 1617.000 ;
      RECT 1201.900 1.400 1202.180 1617.000 ;
      RECT 1204.140 1.400 1204.420 1617.000 ;
      RECT 1206.380 1.400 1206.660 1617.000 ;
      RECT 1208.620 1.400 1208.900 1617.000 ;
      RECT 1210.860 1.400 1211.140 1617.000 ;
      RECT 1213.100 1.400 1213.380 1617.000 ;
      RECT 1215.340 1.400 1215.620 1617.000 ;
      RECT 1217.580 1.400 1217.860 1617.000 ;
      RECT 1219.820 1.400 1220.100 1617.000 ;
      RECT 1222.060 1.400 1222.340 1617.000 ;
      RECT 1224.300 1.400 1224.580 1617.000 ;
      RECT 1226.540 1.400 1226.820 1617.000 ;
      RECT 1228.780 1.400 1229.060 1617.000 ;
      RECT 1231.020 1.400 1231.300 1617.000 ;
      RECT 1233.260 1.400 1233.540 1617.000 ;
      RECT 1235.500 1.400 1235.780 1617.000 ;
      RECT 1237.740 1.400 1238.020 1617.000 ;
      RECT 1239.980 1.400 1240.260 1617.000 ;
      RECT 1242.220 1.400 1242.500 1617.000 ;
      RECT 1244.460 1.400 1244.740 1617.000 ;
      RECT 1246.700 1.400 1246.980 1617.000 ;
      RECT 1248.940 1.400 1249.220 1617.000 ;
      RECT 1251.180 1.400 1251.460 1617.000 ;
      RECT 1253.420 1.400 1253.700 1617.000 ;
      RECT 1255.660 1.400 1255.940 1617.000 ;
      RECT 1257.900 1.400 1258.180 1617.000 ;
      RECT 1260.140 1.400 1260.420 1617.000 ;
      RECT 1262.380 1.400 1262.660 1617.000 ;
      RECT 1264.620 1.400 1264.900 1617.000 ;
      RECT 1266.860 1.400 1267.140 1617.000 ;
      RECT 1269.100 1.400 1269.380 1617.000 ;
      RECT 1271.340 1.400 1271.620 1617.000 ;
      RECT 1273.580 1.400 1273.860 1617.000 ;
      RECT 1275.820 1.400 1276.100 1617.000 ;
      RECT 1278.060 1.400 1278.340 1617.000 ;
      RECT 1280.300 1.400 1280.580 1617.000 ;
      RECT 1282.540 1.400 1282.820 1617.000 ;
      RECT 1284.780 1.400 1285.060 1617.000 ;
      RECT 1287.020 1.400 1287.300 1617.000 ;
      RECT 1289.260 1.400 1289.540 1617.000 ;
      RECT 1291.500 1.400 1291.780 1617.000 ;
      RECT 1293.740 1.400 1294.020 1617.000 ;
      RECT 1295.980 1.400 1296.260 1617.000 ;
      RECT 1298.220 1.400 1298.500 1617.000 ;
      RECT 1300.460 1.400 1300.740 1617.000 ;
      RECT 1302.700 1.400 1302.980 1617.000 ;
      RECT 1304.940 1.400 1305.220 1617.000 ;
      RECT 1307.180 1.400 1307.460 1617.000 ;
      RECT 1309.420 1.400 1309.700 1617.000 ;
      RECT 1311.660 1.400 1311.940 1617.000 ;
      RECT 1313.900 1.400 1314.180 1617.000 ;
      RECT 1316.140 1.400 1316.420 1617.000 ;
      RECT 1318.380 1.400 1318.660 1617.000 ;
      RECT 1320.620 1.400 1320.900 1617.000 ;
      RECT 1322.860 1.400 1323.140 1617.000 ;
      RECT 1325.100 1.400 1325.380 1617.000 ;
      RECT 1327.340 1.400 1327.620 1617.000 ;
      RECT 1329.580 1.400 1329.860 1617.000 ;
      RECT 1331.820 1.400 1332.100 1617.000 ;
      RECT 1334.060 1.400 1334.340 1617.000 ;
      RECT 1336.300 1.400 1336.580 1617.000 ;
      RECT 1338.540 1.400 1338.820 1617.000 ;
      RECT 1340.780 1.400 1341.060 1617.000 ;
      RECT 1343.020 1.400 1343.300 1617.000 ;
      RECT 1345.260 1.400 1345.540 1617.000 ;
      RECT 1347.500 1.400 1347.780 1617.000 ;
      RECT 1349.740 1.400 1350.020 1617.000 ;
      RECT 1351.980 1.400 1352.260 1617.000 ;
      RECT 1354.220 1.400 1354.500 1617.000 ;
      RECT 1356.460 1.400 1356.740 1617.000 ;
      RECT 1358.700 1.400 1358.980 1617.000 ;
      RECT 1360.940 1.400 1361.220 1617.000 ;
      RECT 1363.180 1.400 1363.460 1617.000 ;
      RECT 1365.420 1.400 1365.700 1617.000 ;
      RECT 1367.660 1.400 1367.940 1617.000 ;
      RECT 1369.900 1.400 1370.180 1617.000 ;
      RECT 1372.140 1.400 1372.420 1617.000 ;
      RECT 1374.380 1.400 1374.660 1617.000 ;
      RECT 1376.620 1.400 1376.900 1617.000 ;
      RECT 1378.860 1.400 1379.140 1617.000 ;
      RECT 1381.100 1.400 1381.380 1617.000 ;
      RECT 1383.340 1.400 1383.620 1617.000 ;
      RECT 1385.580 1.400 1385.860 1617.000 ;
      RECT 1387.820 1.400 1388.100 1617.000 ;
      RECT 1390.060 1.400 1390.340 1617.000 ;
      RECT 1392.300 1.400 1392.580 1617.000 ;
      RECT 1394.540 1.400 1394.820 1617.000 ;
      RECT 1396.780 1.400 1397.060 1617.000 ;
      RECT 1399.020 1.400 1399.300 1617.000 ;
      RECT 1401.260 1.400 1401.540 1617.000 ;
      RECT 1403.500 1.400 1403.780 1617.000 ;
      RECT 1405.740 1.400 1406.020 1617.000 ;
      RECT 1407.980 1.400 1408.260 1617.000 ;
      RECT 1410.220 1.400 1410.500 1617.000 ;
      RECT 1412.460 1.400 1412.740 1617.000 ;
      RECT 1414.700 1.400 1414.980 1617.000 ;
      RECT 1416.940 1.400 1417.220 1617.000 ;
      RECT 1419.180 1.400 1419.460 1617.000 ;
      RECT 1421.420 1.400 1421.700 1617.000 ;
      RECT 1423.660 1.400 1423.940 1617.000 ;
      RECT 1425.900 1.400 1426.180 1617.000 ;
      RECT 1428.140 1.400 1428.420 1617.000 ;
      RECT 1430.380 1.400 1430.660 1617.000 ;
      RECT 1432.620 1.400 1432.900 1617.000 ;
      RECT 1434.860 1.400 1435.140 1617.000 ;
      RECT 1437.100 1.400 1437.380 1617.000 ;
      RECT 1439.340 1.400 1439.620 1617.000 ;
      RECT 1441.580 1.400 1441.860 1617.000 ;
      RECT 1443.820 1.400 1444.100 1617.000 ;
      RECT 1446.060 1.400 1446.340 1617.000 ;
      RECT 1448.300 1.400 1448.580 1617.000 ;
      RECT 1450.540 1.400 1450.820 1617.000 ;
      RECT 1452.780 1.400 1453.060 1617.000 ;
      RECT 1455.020 1.400 1455.300 1617.000 ;
      RECT 1457.260 1.400 1457.540 1617.000 ;
      RECT 1459.500 1.400 1459.780 1617.000 ;
      RECT 1461.740 1.400 1462.020 1617.000 ;
      RECT 1463.980 1.400 1464.260 1617.000 ;
      RECT 1466.220 1.400 1466.500 1617.000 ;
      RECT 1468.460 1.400 1468.740 1617.000 ;
      RECT 1470.700 1.400 1470.980 1617.000 ;
      RECT 1472.940 1.400 1473.220 1617.000 ;
      RECT 1475.180 1.400 1475.460 1617.000 ;
      RECT 1477.420 1.400 1477.700 1617.000 ;
      RECT 1479.660 1.400 1479.940 1617.000 ;
      RECT 1481.900 1.400 1482.180 1617.000 ;
      RECT 1484.140 1.400 1484.420 1617.000 ;
      RECT 1486.380 1.400 1486.660 1617.000 ;
      RECT 1488.620 1.400 1488.900 1617.000 ;
      RECT 1490.860 1.400 1491.140 1617.000 ;
      RECT 1493.100 1.400 1493.380 1617.000 ;
      RECT 1495.340 1.400 1495.620 1617.000 ;
      RECT 1497.580 1.400 1497.860 1617.000 ;
      RECT 1499.820 1.400 1500.100 1617.000 ;
      RECT 1502.060 1.400 1502.340 1617.000 ;
      RECT 1504.300 1.400 1504.580 1617.000 ;
      RECT 1506.540 1.400 1506.820 1617.000 ;
      RECT 1508.780 1.400 1509.060 1617.000 ;
      RECT 1511.020 1.400 1511.300 1617.000 ;
      RECT 1513.260 1.400 1513.540 1617.000 ;
      RECT 1515.500 1.400 1515.780 1617.000 ;
      RECT 1517.740 1.400 1518.020 1617.000 ;
      RECT 1519.980 1.400 1520.260 1617.000 ;
      RECT 1522.220 1.400 1522.500 1617.000 ;
      RECT 1524.460 1.400 1524.740 1617.000 ;
      RECT 1526.700 1.400 1526.980 1617.000 ;
      RECT 1528.940 1.400 1529.220 1617.000 ;
      RECT 1531.180 1.400 1531.460 1617.000 ;
      RECT 1533.420 1.400 1533.700 1617.000 ;
      RECT 1535.660 1.400 1535.940 1617.000 ;
      RECT 1537.900 1.400 1538.180 1617.000 ;
      RECT 1540.140 1.400 1540.420 1617.000 ;
      RECT 1542.380 1.400 1542.660 1617.000 ;
      RECT 1544.620 1.400 1544.900 1617.000 ;
      RECT 1546.860 1.400 1547.140 1617.000 ;
      RECT 1549.100 1.400 1549.380 1617.000 ;
      RECT 1551.340 1.400 1551.620 1617.000 ;
      RECT 1553.580 1.400 1553.860 1617.000 ;
      RECT 1555.820 1.400 1556.100 1617.000 ;
      RECT 1558.060 1.400 1558.340 1617.000 ;
      RECT 1560.300 1.400 1560.580 1617.000 ;
      RECT 1562.540 1.400 1562.820 1617.000 ;
      RECT 1564.780 1.400 1565.060 1617.000 ;
      RECT 1567.020 1.400 1567.300 1617.000 ;
      RECT 1569.260 1.400 1569.540 1617.000 ;
      RECT 1571.500 1.400 1571.780 1617.000 ;
      RECT 1573.740 1.400 1574.020 1617.000 ;
      RECT 1575.980 1.400 1576.260 1617.000 ;
      RECT 1578.220 1.400 1578.500 1617.000 ;
      RECT 1580.460 1.400 1580.740 1617.000 ;
      RECT 1582.700 1.400 1582.980 1617.000 ;
      RECT 1584.940 1.400 1585.220 1617.000 ;
      RECT 1587.180 1.400 1587.460 1617.000 ;
      RECT 1589.420 1.400 1589.700 1617.000 ;
      RECT 1591.660 1.400 1591.940 1617.000 ;
      RECT 1593.900 1.400 1594.180 1617.000 ;
      RECT 1596.140 1.400 1596.420 1617.000 ;
      RECT 1598.380 1.400 1598.660 1617.000 ;
      RECT 1600.620 1.400 1600.900 1617.000 ;
      RECT 1602.860 1.400 1603.140 1617.000 ;
      RECT 1605.100 1.400 1605.380 1617.000 ;
      RECT 1607.340 1.400 1607.620 1617.000 ;
      RECT 1609.580 1.400 1609.860 1617.000 ;
      RECT 1611.820 1.400 1612.100 1617.000 ;
      RECT 1614.060 1.400 1614.340 1617.000 ;
      RECT 1616.300 1.400 1616.580 1617.000 ;
      RECT 1618.540 1.400 1618.820 1617.000 ;
      RECT 1620.780 1.400 1621.060 1617.000 ;
      RECT 1623.020 1.400 1623.300 1617.000 ;
      RECT 1625.260 1.400 1625.540 1617.000 ;
      RECT 1627.500 1.400 1627.780 1617.000 ;
      RECT 1629.740 1.400 1630.020 1617.000 ;
      RECT 1631.980 1.400 1632.260 1617.000 ;
      RECT 1634.220 1.400 1634.500 1617.000 ;
      RECT 1636.460 1.400 1636.740 1617.000 ;
      RECT 1638.700 1.400 1638.980 1617.000 ;
      RECT 1640.940 1.400 1641.220 1617.000 ;
      RECT 1643.180 1.400 1643.460 1617.000 ;
      RECT 1645.420 1.400 1645.700 1617.000 ;
      RECT 1647.660 1.400 1647.940 1617.000 ;
      RECT 1649.900 1.400 1650.180 1617.000 ;
      RECT 1652.140 1.400 1652.420 1617.000 ;
      RECT 1654.380 1.400 1654.660 1617.000 ;
      RECT 1656.620 1.400 1656.900 1617.000 ;
      RECT 1658.860 1.400 1659.140 1617.000 ;
      RECT 1661.100 1.400 1661.380 1617.000 ;
      RECT 1663.340 1.400 1663.620 1617.000 ;
      RECT 1665.580 1.400 1665.860 1617.000 ;
      RECT 1667.820 1.400 1668.100 1617.000 ;
      RECT 1670.060 1.400 1670.340 1617.000 ;
      RECT 1672.300 1.400 1672.580 1617.000 ;
      RECT 1674.540 1.400 1674.820 1617.000 ;
      RECT 1676.780 1.400 1677.060 1617.000 ;
      RECT 1679.020 1.400 1679.300 1617.000 ;
      RECT 1681.260 1.400 1681.540 1617.000 ;
      RECT 1683.500 1.400 1683.780 1617.000 ;
      RECT 1685.740 1.400 1686.020 1617.000 ;
      RECT 1687.980 1.400 1688.260 1617.000 ;
      RECT 1690.220 1.400 1690.500 1617.000 ;
      RECT 1692.460 1.400 1692.740 1617.000 ;
      RECT 1694.700 1.400 1694.980 1617.000 ;
      RECT 1696.940 1.400 1697.220 1617.000 ;
      RECT 1699.180 1.400 1699.460 1617.000 ;
      RECT 1701.420 1.400 1701.700 1617.000 ;
      RECT 1703.660 1.400 1703.940 1617.000 ;
      RECT 1705.900 1.400 1706.180 1617.000 ;
      RECT 1708.140 1.400 1708.420 1617.000 ;
      RECT 1710.380 1.400 1710.660 1617.000 ;
      RECT 1712.620 1.400 1712.900 1617.000 ;
      RECT 1714.860 1.400 1715.140 1617.000 ;
      RECT 1717.100 1.400 1717.380 1617.000 ;
      RECT 1719.340 1.400 1719.620 1617.000 ;
      RECT 1721.580 1.400 1721.860 1617.000 ;
      RECT 1723.820 1.400 1724.100 1617.000 ;
      RECT 1726.060 1.400 1726.340 1617.000 ;
      RECT 1728.300 1.400 1728.580 1617.000 ;
      RECT 1730.540 1.400 1730.820 1617.000 ;
      RECT 1732.780 1.400 1733.060 1617.000 ;
      RECT 1735.020 1.400 1735.300 1617.000 ;
      RECT 1737.260 1.400 1737.540 1617.000 ;
      RECT 1739.500 1.400 1739.780 1617.000 ;
      RECT 1741.740 1.400 1742.020 1617.000 ;
      RECT 1743.980 1.400 1744.260 1617.000 ;
      RECT 1746.220 1.400 1746.500 1617.000 ;
      RECT 1748.460 1.400 1748.740 1617.000 ;
      RECT 1750.700 1.400 1750.980 1617.000 ;
      RECT 1752.940 1.400 1753.220 1617.000 ;
      RECT 1755.180 1.400 1755.460 1617.000 ;
      RECT 1757.420 1.400 1757.700 1617.000 ;
      RECT 1759.660 1.400 1759.940 1617.000 ;
      RECT 1761.900 1.400 1762.180 1617.000 ;
      RECT 1764.140 1.400 1764.420 1617.000 ;
      RECT 1766.380 1.400 1766.660 1617.000 ;
      RECT 1768.620 1.400 1768.900 1617.000 ;
      RECT 1770.860 1.400 1771.140 1617.000 ;
      RECT 1773.100 1.400 1773.380 1617.000 ;
      RECT 1775.340 1.400 1775.620 1617.000 ;
      RECT 1777.580 1.400 1777.860 1617.000 ;
      RECT 1779.820 1.400 1780.100 1617.000 ;
      RECT 1782.060 1.400 1782.340 1617.000 ;
      RECT 1784.300 1.400 1784.580 1617.000 ;
      RECT 1786.540 1.400 1786.820 1617.000 ;
      RECT 1788.780 1.400 1789.060 1617.000 ;
      RECT 1791.020 1.400 1791.300 1617.000 ;
      RECT 1793.260 1.400 1793.540 1617.000 ;
      RECT 1795.500 1.400 1795.780 1617.000 ;
      RECT 1797.740 1.400 1798.020 1617.000 ;
      RECT 1799.980 1.400 1800.260 1617.000 ;
      RECT 1802.220 1.400 1802.500 1617.000 ;
      RECT 1804.460 1.400 1804.740 1617.000 ;
      RECT 1806.700 1.400 1806.980 1617.000 ;
      RECT 1808.940 1.400 1809.220 1617.000 ;
      RECT 1811.180 1.400 1811.460 1617.000 ;
      RECT 1813.420 1.400 1813.700 1617.000 ;
      RECT 1815.660 1.400 1815.940 1617.000 ;
      RECT 1817.900 1.400 1818.180 1617.000 ;
      RECT 1820.140 1.400 1820.420 1617.000 ;
      RECT 1822.380 1.400 1822.660 1617.000 ;
      RECT 1824.620 1.400 1824.900 1617.000 ;
      RECT 1826.860 1.400 1827.140 1617.000 ;
      RECT 1829.100 1.400 1829.380 1617.000 ;
      RECT 1831.340 1.400 1831.620 1617.000 ;
      RECT 1833.580 1.400 1833.860 1617.000 ;
      RECT 1835.820 1.400 1836.100 1617.000 ;
      RECT 1838.060 1.400 1838.340 1617.000 ;
      RECT 1840.300 1.400 1840.580 1617.000 ;
      RECT 1842.540 1.400 1842.820 1617.000 ;
      RECT 1844.780 1.400 1845.060 1617.000 ;
      RECT 1847.020 1.400 1847.300 1617.000 ;
      RECT 1849.260 1.400 1849.540 1617.000 ;
      RECT 1851.500 1.400 1851.780 1617.000 ;
      RECT 1853.740 1.400 1854.020 1617.000 ;
      RECT 1855.980 1.400 1856.260 1617.000 ;
      RECT 1858.220 1.400 1858.500 1617.000 ;
      RECT 1860.460 1.400 1860.740 1617.000 ;
      RECT 1862.700 1.400 1862.980 1617.000 ;
      RECT 1864.940 1.400 1865.220 1617.000 ;
      RECT 1867.180 1.400 1867.460 1617.000 ;
      RECT 1869.420 1.400 1869.700 1617.000 ;
      RECT 1871.660 1.400 1871.940 1617.000 ;
      RECT 1873.900 1.400 1874.180 1617.000 ;
      RECT 1876.140 1.400 1876.420 1617.000 ;
      RECT 1878.380 1.400 1878.660 1617.000 ;
      RECT 1880.620 1.400 1880.900 1617.000 ;
      RECT 1882.860 1.400 1883.140 1617.000 ;
      RECT 1885.100 1.400 1885.380 1617.000 ;
      RECT 1887.340 1.400 1887.620 1617.000 ;
      RECT 1889.580 1.400 1889.860 1617.000 ;
      RECT 1891.820 1.400 1892.100 1617.000 ;
      RECT 1894.060 1.400 1894.340 1617.000 ;
      RECT 1896.300 1.400 1896.580 1617.000 ;
      RECT 1898.540 1.400 1898.820 1617.000 ;
      RECT 1900.780 1.400 1901.060 1617.000 ;
      RECT 1903.020 1.400 1903.300 1617.000 ;
      RECT 1905.260 1.400 1905.540 1617.000 ;
      RECT 1907.500 1.400 1907.780 1617.000 ;
      RECT 1909.740 1.400 1910.020 1617.000 ;
      RECT 1911.980 1.400 1912.260 1617.000 ;
      RECT 1914.220 1.400 1914.500 1617.000 ;
      RECT 1916.460 1.400 1916.740 1617.000 ;
      RECT 1918.700 1.400 1918.980 1617.000 ;
      RECT 1920.940 1.400 1921.220 1617.000 ;
      RECT 1923.180 1.400 1923.460 1617.000 ;
      RECT 1925.420 1.400 1925.700 1617.000 ;
      RECT 1927.660 1.400 1927.940 1617.000 ;
      RECT 1929.900 1.400 1930.180 1617.000 ;
      RECT 1932.140 1.400 1932.420 1617.000 ;
      RECT 1934.380 1.400 1934.660 1617.000 ;
      RECT 1936.620 1.400 1936.900 1617.000 ;
      RECT 1938.860 1.400 1939.140 1617.000 ;
      RECT 1941.100 1.400 1941.380 1617.000 ;
      RECT 1943.340 1.400 1943.620 1617.000 ;
      RECT 1945.580 1.400 1945.860 1617.000 ;
      RECT 1947.820 1.400 1948.100 1617.000 ;
      RECT 1950.060 1.400 1950.340 1617.000 ;
      RECT 1952.300 1.400 1952.580 1617.000 ;
      RECT 1954.540 1.400 1954.820 1617.000 ;
      RECT 1956.780 1.400 1957.060 1617.000 ;
      RECT 1959.020 1.400 1959.300 1617.000 ;
      RECT 1961.260 1.400 1961.540 1617.000 ;
      RECT 1963.500 1.400 1963.780 1617.000 ;
      RECT 1965.740 1.400 1966.020 1617.000 ;
      RECT 1967.980 1.400 1968.260 1617.000 ;
      RECT 1970.220 1.400 1970.500 1617.000 ;
      RECT 1972.460 1.400 1972.740 1617.000 ;
      RECT 1974.700 1.400 1974.980 1617.000 ;
      RECT 1976.940 1.400 1977.220 1617.000 ;
      RECT 1979.180 1.400 1979.460 1617.000 ;
      RECT 1981.420 1.400 1981.700 1617.000 ;
      RECT 1983.660 1.400 1983.940 1617.000 ;
      RECT 1985.900 1.400 1986.180 1617.000 ;
      RECT 1988.140 1.400 1988.420 1617.000 ;
      RECT 1990.380 1.400 1990.660 1617.000 ;
      RECT 1992.620 1.400 1992.900 1617.000 ;
      RECT 1994.860 1.400 1995.140 1617.000 ;
      RECT 1997.100 1.400 1997.380 1617.000 ;
      RECT 1999.340 1.400 1999.620 1617.000 ;
      RECT 2001.580 1.400 2001.860 1617.000 ;
      RECT 2003.820 1.400 2004.100 1617.000 ;
      RECT 2006.060 1.400 2006.340 1617.000 ;
      RECT 2008.300 1.400 2008.580 1617.000 ;
      RECT 2010.540 1.400 2010.820 1617.000 ;
      RECT 2012.780 1.400 2013.060 1617.000 ;
      RECT 2015.020 1.400 2015.300 1617.000 ;
      RECT 2017.260 1.400 2017.540 1617.000 ;
      RECT 2019.500 1.400 2019.780 1617.000 ;
      RECT 2021.740 1.400 2022.020 1617.000 ;
      RECT 2023.980 1.400 2024.260 1617.000 ;
      RECT 2026.220 1.400 2026.500 1617.000 ;
      RECT 2028.460 1.400 2028.740 1617.000 ;
      RECT 2030.700 1.400 2030.980 1617.000 ;
      RECT 2032.940 1.400 2033.220 1617.000 ;
      RECT 2035.180 1.400 2035.460 1617.000 ;
      RECT 2037.420 1.400 2037.700 1617.000 ;
      RECT 2039.660 1.400 2039.940 1617.000 ;
      RECT 2041.900 1.400 2042.180 1617.000 ;
      RECT 2044.140 1.400 2044.420 1617.000 ;
      RECT 2046.380 1.400 2046.660 1617.000 ;
      RECT 2048.620 1.400 2048.900 1617.000 ;
      RECT 2050.860 1.400 2051.140 1617.000 ;
      RECT 2053.100 1.400 2053.380 1617.000 ;
      RECT 2055.340 1.400 2055.620 1617.000 ;
      RECT 2057.580 1.400 2057.860 1617.000 ;
      RECT 2059.820 1.400 2060.100 1617.000 ;
      RECT 2062.060 1.400 2062.340 1617.000 ;
      RECT 2064.300 1.400 2064.580 1617.000 ;
      RECT 2066.540 1.400 2066.820 1617.000 ;
      RECT 2068.780 1.400 2069.060 1617.000 ;
      RECT 2071.020 1.400 2071.300 1617.000 ;
      RECT 2073.260 1.400 2073.540 1617.000 ;
      RECT 2075.500 1.400 2075.780 1617.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 1617.000 ;
      RECT 4.620 1.400 4.900 1617.000 ;
      RECT 6.860 1.400 7.140 1617.000 ;
      RECT 9.100 1.400 9.380 1617.000 ;
      RECT 11.340 1.400 11.620 1617.000 ;
      RECT 13.580 1.400 13.860 1617.000 ;
      RECT 15.820 1.400 16.100 1617.000 ;
      RECT 18.060 1.400 18.340 1617.000 ;
      RECT 20.300 1.400 20.580 1617.000 ;
      RECT 22.540 1.400 22.820 1617.000 ;
      RECT 24.780 1.400 25.060 1617.000 ;
      RECT 27.020 1.400 27.300 1617.000 ;
      RECT 29.260 1.400 29.540 1617.000 ;
      RECT 31.500 1.400 31.780 1617.000 ;
      RECT 33.740 1.400 34.020 1617.000 ;
      RECT 35.980 1.400 36.260 1617.000 ;
      RECT 38.220 1.400 38.500 1617.000 ;
      RECT 40.460 1.400 40.740 1617.000 ;
      RECT 42.700 1.400 42.980 1617.000 ;
      RECT 44.940 1.400 45.220 1617.000 ;
      RECT 47.180 1.400 47.460 1617.000 ;
      RECT 49.420 1.400 49.700 1617.000 ;
      RECT 51.660 1.400 51.940 1617.000 ;
      RECT 53.900 1.400 54.180 1617.000 ;
      RECT 56.140 1.400 56.420 1617.000 ;
      RECT 58.380 1.400 58.660 1617.000 ;
      RECT 60.620 1.400 60.900 1617.000 ;
      RECT 62.860 1.400 63.140 1617.000 ;
      RECT 65.100 1.400 65.380 1617.000 ;
      RECT 67.340 1.400 67.620 1617.000 ;
      RECT 69.580 1.400 69.860 1617.000 ;
      RECT 71.820 1.400 72.100 1617.000 ;
      RECT 74.060 1.400 74.340 1617.000 ;
      RECT 76.300 1.400 76.580 1617.000 ;
      RECT 78.540 1.400 78.820 1617.000 ;
      RECT 80.780 1.400 81.060 1617.000 ;
      RECT 83.020 1.400 83.300 1617.000 ;
      RECT 85.260 1.400 85.540 1617.000 ;
      RECT 87.500 1.400 87.780 1617.000 ;
      RECT 89.740 1.400 90.020 1617.000 ;
      RECT 91.980 1.400 92.260 1617.000 ;
      RECT 94.220 1.400 94.500 1617.000 ;
      RECT 96.460 1.400 96.740 1617.000 ;
      RECT 98.700 1.400 98.980 1617.000 ;
      RECT 100.940 1.400 101.220 1617.000 ;
      RECT 103.180 1.400 103.460 1617.000 ;
      RECT 105.420 1.400 105.700 1617.000 ;
      RECT 107.660 1.400 107.940 1617.000 ;
      RECT 109.900 1.400 110.180 1617.000 ;
      RECT 112.140 1.400 112.420 1617.000 ;
      RECT 114.380 1.400 114.660 1617.000 ;
      RECT 116.620 1.400 116.900 1617.000 ;
      RECT 118.860 1.400 119.140 1617.000 ;
      RECT 121.100 1.400 121.380 1617.000 ;
      RECT 123.340 1.400 123.620 1617.000 ;
      RECT 125.580 1.400 125.860 1617.000 ;
      RECT 127.820 1.400 128.100 1617.000 ;
      RECT 130.060 1.400 130.340 1617.000 ;
      RECT 132.300 1.400 132.580 1617.000 ;
      RECT 134.540 1.400 134.820 1617.000 ;
      RECT 136.780 1.400 137.060 1617.000 ;
      RECT 139.020 1.400 139.300 1617.000 ;
      RECT 141.260 1.400 141.540 1617.000 ;
      RECT 143.500 1.400 143.780 1617.000 ;
      RECT 145.740 1.400 146.020 1617.000 ;
      RECT 147.980 1.400 148.260 1617.000 ;
      RECT 150.220 1.400 150.500 1617.000 ;
      RECT 152.460 1.400 152.740 1617.000 ;
      RECT 154.700 1.400 154.980 1617.000 ;
      RECT 156.940 1.400 157.220 1617.000 ;
      RECT 159.180 1.400 159.460 1617.000 ;
      RECT 161.420 1.400 161.700 1617.000 ;
      RECT 163.660 1.400 163.940 1617.000 ;
      RECT 165.900 1.400 166.180 1617.000 ;
      RECT 168.140 1.400 168.420 1617.000 ;
      RECT 170.380 1.400 170.660 1617.000 ;
      RECT 172.620 1.400 172.900 1617.000 ;
      RECT 174.860 1.400 175.140 1617.000 ;
      RECT 177.100 1.400 177.380 1617.000 ;
      RECT 179.340 1.400 179.620 1617.000 ;
      RECT 181.580 1.400 181.860 1617.000 ;
      RECT 183.820 1.400 184.100 1617.000 ;
      RECT 186.060 1.400 186.340 1617.000 ;
      RECT 188.300 1.400 188.580 1617.000 ;
      RECT 190.540 1.400 190.820 1617.000 ;
      RECT 192.780 1.400 193.060 1617.000 ;
      RECT 195.020 1.400 195.300 1617.000 ;
      RECT 197.260 1.400 197.540 1617.000 ;
      RECT 199.500 1.400 199.780 1617.000 ;
      RECT 201.740 1.400 202.020 1617.000 ;
      RECT 203.980 1.400 204.260 1617.000 ;
      RECT 206.220 1.400 206.500 1617.000 ;
      RECT 208.460 1.400 208.740 1617.000 ;
      RECT 210.700 1.400 210.980 1617.000 ;
      RECT 212.940 1.400 213.220 1617.000 ;
      RECT 215.180 1.400 215.460 1617.000 ;
      RECT 217.420 1.400 217.700 1617.000 ;
      RECT 219.660 1.400 219.940 1617.000 ;
      RECT 221.900 1.400 222.180 1617.000 ;
      RECT 224.140 1.400 224.420 1617.000 ;
      RECT 226.380 1.400 226.660 1617.000 ;
      RECT 228.620 1.400 228.900 1617.000 ;
      RECT 230.860 1.400 231.140 1617.000 ;
      RECT 233.100 1.400 233.380 1617.000 ;
      RECT 235.340 1.400 235.620 1617.000 ;
      RECT 237.580 1.400 237.860 1617.000 ;
      RECT 239.820 1.400 240.100 1617.000 ;
      RECT 242.060 1.400 242.340 1617.000 ;
      RECT 244.300 1.400 244.580 1617.000 ;
      RECT 246.540 1.400 246.820 1617.000 ;
      RECT 248.780 1.400 249.060 1617.000 ;
      RECT 251.020 1.400 251.300 1617.000 ;
      RECT 253.260 1.400 253.540 1617.000 ;
      RECT 255.500 1.400 255.780 1617.000 ;
      RECT 257.740 1.400 258.020 1617.000 ;
      RECT 259.980 1.400 260.260 1617.000 ;
      RECT 262.220 1.400 262.500 1617.000 ;
      RECT 264.460 1.400 264.740 1617.000 ;
      RECT 266.700 1.400 266.980 1617.000 ;
      RECT 268.940 1.400 269.220 1617.000 ;
      RECT 271.180 1.400 271.460 1617.000 ;
      RECT 273.420 1.400 273.700 1617.000 ;
      RECT 275.660 1.400 275.940 1617.000 ;
      RECT 277.900 1.400 278.180 1617.000 ;
      RECT 280.140 1.400 280.420 1617.000 ;
      RECT 282.380 1.400 282.660 1617.000 ;
      RECT 284.620 1.400 284.900 1617.000 ;
      RECT 286.860 1.400 287.140 1617.000 ;
      RECT 289.100 1.400 289.380 1617.000 ;
      RECT 291.340 1.400 291.620 1617.000 ;
      RECT 293.580 1.400 293.860 1617.000 ;
      RECT 295.820 1.400 296.100 1617.000 ;
      RECT 298.060 1.400 298.340 1617.000 ;
      RECT 300.300 1.400 300.580 1617.000 ;
      RECT 302.540 1.400 302.820 1617.000 ;
      RECT 304.780 1.400 305.060 1617.000 ;
      RECT 307.020 1.400 307.300 1617.000 ;
      RECT 309.260 1.400 309.540 1617.000 ;
      RECT 311.500 1.400 311.780 1617.000 ;
      RECT 313.740 1.400 314.020 1617.000 ;
      RECT 315.980 1.400 316.260 1617.000 ;
      RECT 318.220 1.400 318.500 1617.000 ;
      RECT 320.460 1.400 320.740 1617.000 ;
      RECT 322.700 1.400 322.980 1617.000 ;
      RECT 324.940 1.400 325.220 1617.000 ;
      RECT 327.180 1.400 327.460 1617.000 ;
      RECT 329.420 1.400 329.700 1617.000 ;
      RECT 331.660 1.400 331.940 1617.000 ;
      RECT 333.900 1.400 334.180 1617.000 ;
      RECT 336.140 1.400 336.420 1617.000 ;
      RECT 338.380 1.400 338.660 1617.000 ;
      RECT 340.620 1.400 340.900 1617.000 ;
      RECT 342.860 1.400 343.140 1617.000 ;
      RECT 345.100 1.400 345.380 1617.000 ;
      RECT 347.340 1.400 347.620 1617.000 ;
      RECT 349.580 1.400 349.860 1617.000 ;
      RECT 351.820 1.400 352.100 1617.000 ;
      RECT 354.060 1.400 354.340 1617.000 ;
      RECT 356.300 1.400 356.580 1617.000 ;
      RECT 358.540 1.400 358.820 1617.000 ;
      RECT 360.780 1.400 361.060 1617.000 ;
      RECT 363.020 1.400 363.300 1617.000 ;
      RECT 365.260 1.400 365.540 1617.000 ;
      RECT 367.500 1.400 367.780 1617.000 ;
      RECT 369.740 1.400 370.020 1617.000 ;
      RECT 371.980 1.400 372.260 1617.000 ;
      RECT 374.220 1.400 374.500 1617.000 ;
      RECT 376.460 1.400 376.740 1617.000 ;
      RECT 378.700 1.400 378.980 1617.000 ;
      RECT 380.940 1.400 381.220 1617.000 ;
      RECT 383.180 1.400 383.460 1617.000 ;
      RECT 385.420 1.400 385.700 1617.000 ;
      RECT 387.660 1.400 387.940 1617.000 ;
      RECT 389.900 1.400 390.180 1617.000 ;
      RECT 392.140 1.400 392.420 1617.000 ;
      RECT 394.380 1.400 394.660 1617.000 ;
      RECT 396.620 1.400 396.900 1617.000 ;
      RECT 398.860 1.400 399.140 1617.000 ;
      RECT 401.100 1.400 401.380 1617.000 ;
      RECT 403.340 1.400 403.620 1617.000 ;
      RECT 405.580 1.400 405.860 1617.000 ;
      RECT 407.820 1.400 408.100 1617.000 ;
      RECT 410.060 1.400 410.340 1617.000 ;
      RECT 412.300 1.400 412.580 1617.000 ;
      RECT 414.540 1.400 414.820 1617.000 ;
      RECT 416.780 1.400 417.060 1617.000 ;
      RECT 419.020 1.400 419.300 1617.000 ;
      RECT 421.260 1.400 421.540 1617.000 ;
      RECT 423.500 1.400 423.780 1617.000 ;
      RECT 425.740 1.400 426.020 1617.000 ;
      RECT 427.980 1.400 428.260 1617.000 ;
      RECT 430.220 1.400 430.500 1617.000 ;
      RECT 432.460 1.400 432.740 1617.000 ;
      RECT 434.700 1.400 434.980 1617.000 ;
      RECT 436.940 1.400 437.220 1617.000 ;
      RECT 439.180 1.400 439.460 1617.000 ;
      RECT 441.420 1.400 441.700 1617.000 ;
      RECT 443.660 1.400 443.940 1617.000 ;
      RECT 445.900 1.400 446.180 1617.000 ;
      RECT 448.140 1.400 448.420 1617.000 ;
      RECT 450.380 1.400 450.660 1617.000 ;
      RECT 452.620 1.400 452.900 1617.000 ;
      RECT 454.860 1.400 455.140 1617.000 ;
      RECT 457.100 1.400 457.380 1617.000 ;
      RECT 459.340 1.400 459.620 1617.000 ;
      RECT 461.580 1.400 461.860 1617.000 ;
      RECT 463.820 1.400 464.100 1617.000 ;
      RECT 466.060 1.400 466.340 1617.000 ;
      RECT 468.300 1.400 468.580 1617.000 ;
      RECT 470.540 1.400 470.820 1617.000 ;
      RECT 472.780 1.400 473.060 1617.000 ;
      RECT 475.020 1.400 475.300 1617.000 ;
      RECT 477.260 1.400 477.540 1617.000 ;
      RECT 479.500 1.400 479.780 1617.000 ;
      RECT 481.740 1.400 482.020 1617.000 ;
      RECT 483.980 1.400 484.260 1617.000 ;
      RECT 486.220 1.400 486.500 1617.000 ;
      RECT 488.460 1.400 488.740 1617.000 ;
      RECT 490.700 1.400 490.980 1617.000 ;
      RECT 492.940 1.400 493.220 1617.000 ;
      RECT 495.180 1.400 495.460 1617.000 ;
      RECT 497.420 1.400 497.700 1617.000 ;
      RECT 499.660 1.400 499.940 1617.000 ;
      RECT 501.900 1.400 502.180 1617.000 ;
      RECT 504.140 1.400 504.420 1617.000 ;
      RECT 506.380 1.400 506.660 1617.000 ;
      RECT 508.620 1.400 508.900 1617.000 ;
      RECT 510.860 1.400 511.140 1617.000 ;
      RECT 513.100 1.400 513.380 1617.000 ;
      RECT 515.340 1.400 515.620 1617.000 ;
      RECT 517.580 1.400 517.860 1617.000 ;
      RECT 519.820 1.400 520.100 1617.000 ;
      RECT 522.060 1.400 522.340 1617.000 ;
      RECT 524.300 1.400 524.580 1617.000 ;
      RECT 526.540 1.400 526.820 1617.000 ;
      RECT 528.780 1.400 529.060 1617.000 ;
      RECT 531.020 1.400 531.300 1617.000 ;
      RECT 533.260 1.400 533.540 1617.000 ;
      RECT 535.500 1.400 535.780 1617.000 ;
      RECT 537.740 1.400 538.020 1617.000 ;
      RECT 539.980 1.400 540.260 1617.000 ;
      RECT 542.220 1.400 542.500 1617.000 ;
      RECT 544.460 1.400 544.740 1617.000 ;
      RECT 546.700 1.400 546.980 1617.000 ;
      RECT 548.940 1.400 549.220 1617.000 ;
      RECT 551.180 1.400 551.460 1617.000 ;
      RECT 553.420 1.400 553.700 1617.000 ;
      RECT 555.660 1.400 555.940 1617.000 ;
      RECT 557.900 1.400 558.180 1617.000 ;
      RECT 560.140 1.400 560.420 1617.000 ;
      RECT 562.380 1.400 562.660 1617.000 ;
      RECT 564.620 1.400 564.900 1617.000 ;
      RECT 566.860 1.400 567.140 1617.000 ;
      RECT 569.100 1.400 569.380 1617.000 ;
      RECT 571.340 1.400 571.620 1617.000 ;
      RECT 573.580 1.400 573.860 1617.000 ;
      RECT 575.820 1.400 576.100 1617.000 ;
      RECT 578.060 1.400 578.340 1617.000 ;
      RECT 580.300 1.400 580.580 1617.000 ;
      RECT 582.540 1.400 582.820 1617.000 ;
      RECT 584.780 1.400 585.060 1617.000 ;
      RECT 587.020 1.400 587.300 1617.000 ;
      RECT 589.260 1.400 589.540 1617.000 ;
      RECT 591.500 1.400 591.780 1617.000 ;
      RECT 593.740 1.400 594.020 1617.000 ;
      RECT 595.980 1.400 596.260 1617.000 ;
      RECT 598.220 1.400 598.500 1617.000 ;
      RECT 600.460 1.400 600.740 1617.000 ;
      RECT 602.700 1.400 602.980 1617.000 ;
      RECT 604.940 1.400 605.220 1617.000 ;
      RECT 607.180 1.400 607.460 1617.000 ;
      RECT 609.420 1.400 609.700 1617.000 ;
      RECT 611.660 1.400 611.940 1617.000 ;
      RECT 613.900 1.400 614.180 1617.000 ;
      RECT 616.140 1.400 616.420 1617.000 ;
      RECT 618.380 1.400 618.660 1617.000 ;
      RECT 620.620 1.400 620.900 1617.000 ;
      RECT 622.860 1.400 623.140 1617.000 ;
      RECT 625.100 1.400 625.380 1617.000 ;
      RECT 627.340 1.400 627.620 1617.000 ;
      RECT 629.580 1.400 629.860 1617.000 ;
      RECT 631.820 1.400 632.100 1617.000 ;
      RECT 634.060 1.400 634.340 1617.000 ;
      RECT 636.300 1.400 636.580 1617.000 ;
      RECT 638.540 1.400 638.820 1617.000 ;
      RECT 640.780 1.400 641.060 1617.000 ;
      RECT 643.020 1.400 643.300 1617.000 ;
      RECT 645.260 1.400 645.540 1617.000 ;
      RECT 647.500 1.400 647.780 1617.000 ;
      RECT 649.740 1.400 650.020 1617.000 ;
      RECT 651.980 1.400 652.260 1617.000 ;
      RECT 654.220 1.400 654.500 1617.000 ;
      RECT 656.460 1.400 656.740 1617.000 ;
      RECT 658.700 1.400 658.980 1617.000 ;
      RECT 660.940 1.400 661.220 1617.000 ;
      RECT 663.180 1.400 663.460 1617.000 ;
      RECT 665.420 1.400 665.700 1617.000 ;
      RECT 667.660 1.400 667.940 1617.000 ;
      RECT 669.900 1.400 670.180 1617.000 ;
      RECT 672.140 1.400 672.420 1617.000 ;
      RECT 674.380 1.400 674.660 1617.000 ;
      RECT 676.620 1.400 676.900 1617.000 ;
      RECT 678.860 1.400 679.140 1617.000 ;
      RECT 681.100 1.400 681.380 1617.000 ;
      RECT 683.340 1.400 683.620 1617.000 ;
      RECT 685.580 1.400 685.860 1617.000 ;
      RECT 687.820 1.400 688.100 1617.000 ;
      RECT 690.060 1.400 690.340 1617.000 ;
      RECT 692.300 1.400 692.580 1617.000 ;
      RECT 694.540 1.400 694.820 1617.000 ;
      RECT 696.780 1.400 697.060 1617.000 ;
      RECT 699.020 1.400 699.300 1617.000 ;
      RECT 701.260 1.400 701.540 1617.000 ;
      RECT 703.500 1.400 703.780 1617.000 ;
      RECT 705.740 1.400 706.020 1617.000 ;
      RECT 707.980 1.400 708.260 1617.000 ;
      RECT 710.220 1.400 710.500 1617.000 ;
      RECT 712.460 1.400 712.740 1617.000 ;
      RECT 714.700 1.400 714.980 1617.000 ;
      RECT 716.940 1.400 717.220 1617.000 ;
      RECT 719.180 1.400 719.460 1617.000 ;
      RECT 721.420 1.400 721.700 1617.000 ;
      RECT 723.660 1.400 723.940 1617.000 ;
      RECT 725.900 1.400 726.180 1617.000 ;
      RECT 728.140 1.400 728.420 1617.000 ;
      RECT 730.380 1.400 730.660 1617.000 ;
      RECT 732.620 1.400 732.900 1617.000 ;
      RECT 734.860 1.400 735.140 1617.000 ;
      RECT 737.100 1.400 737.380 1617.000 ;
      RECT 739.340 1.400 739.620 1617.000 ;
      RECT 741.580 1.400 741.860 1617.000 ;
      RECT 743.820 1.400 744.100 1617.000 ;
      RECT 746.060 1.400 746.340 1617.000 ;
      RECT 748.300 1.400 748.580 1617.000 ;
      RECT 750.540 1.400 750.820 1617.000 ;
      RECT 752.780 1.400 753.060 1617.000 ;
      RECT 755.020 1.400 755.300 1617.000 ;
      RECT 757.260 1.400 757.540 1617.000 ;
      RECT 759.500 1.400 759.780 1617.000 ;
      RECT 761.740 1.400 762.020 1617.000 ;
      RECT 763.980 1.400 764.260 1617.000 ;
      RECT 766.220 1.400 766.500 1617.000 ;
      RECT 768.460 1.400 768.740 1617.000 ;
      RECT 770.700 1.400 770.980 1617.000 ;
      RECT 772.940 1.400 773.220 1617.000 ;
      RECT 775.180 1.400 775.460 1617.000 ;
      RECT 777.420 1.400 777.700 1617.000 ;
      RECT 779.660 1.400 779.940 1617.000 ;
      RECT 781.900 1.400 782.180 1617.000 ;
      RECT 784.140 1.400 784.420 1617.000 ;
      RECT 786.380 1.400 786.660 1617.000 ;
      RECT 788.620 1.400 788.900 1617.000 ;
      RECT 790.860 1.400 791.140 1617.000 ;
      RECT 793.100 1.400 793.380 1617.000 ;
      RECT 795.340 1.400 795.620 1617.000 ;
      RECT 797.580 1.400 797.860 1617.000 ;
      RECT 799.820 1.400 800.100 1617.000 ;
      RECT 802.060 1.400 802.340 1617.000 ;
      RECT 804.300 1.400 804.580 1617.000 ;
      RECT 806.540 1.400 806.820 1617.000 ;
      RECT 808.780 1.400 809.060 1617.000 ;
      RECT 811.020 1.400 811.300 1617.000 ;
      RECT 813.260 1.400 813.540 1617.000 ;
      RECT 815.500 1.400 815.780 1617.000 ;
      RECT 817.740 1.400 818.020 1617.000 ;
      RECT 819.980 1.400 820.260 1617.000 ;
      RECT 822.220 1.400 822.500 1617.000 ;
      RECT 824.460 1.400 824.740 1617.000 ;
      RECT 826.700 1.400 826.980 1617.000 ;
      RECT 828.940 1.400 829.220 1617.000 ;
      RECT 831.180 1.400 831.460 1617.000 ;
      RECT 833.420 1.400 833.700 1617.000 ;
      RECT 835.660 1.400 835.940 1617.000 ;
      RECT 837.900 1.400 838.180 1617.000 ;
      RECT 840.140 1.400 840.420 1617.000 ;
      RECT 842.380 1.400 842.660 1617.000 ;
      RECT 844.620 1.400 844.900 1617.000 ;
      RECT 846.860 1.400 847.140 1617.000 ;
      RECT 849.100 1.400 849.380 1617.000 ;
      RECT 851.340 1.400 851.620 1617.000 ;
      RECT 853.580 1.400 853.860 1617.000 ;
      RECT 855.820 1.400 856.100 1617.000 ;
      RECT 858.060 1.400 858.340 1617.000 ;
      RECT 860.300 1.400 860.580 1617.000 ;
      RECT 862.540 1.400 862.820 1617.000 ;
      RECT 864.780 1.400 865.060 1617.000 ;
      RECT 867.020 1.400 867.300 1617.000 ;
      RECT 869.260 1.400 869.540 1617.000 ;
      RECT 871.500 1.400 871.780 1617.000 ;
      RECT 873.740 1.400 874.020 1617.000 ;
      RECT 875.980 1.400 876.260 1617.000 ;
      RECT 878.220 1.400 878.500 1617.000 ;
      RECT 880.460 1.400 880.740 1617.000 ;
      RECT 882.700 1.400 882.980 1617.000 ;
      RECT 884.940 1.400 885.220 1617.000 ;
      RECT 887.180 1.400 887.460 1617.000 ;
      RECT 889.420 1.400 889.700 1617.000 ;
      RECT 891.660 1.400 891.940 1617.000 ;
      RECT 893.900 1.400 894.180 1617.000 ;
      RECT 896.140 1.400 896.420 1617.000 ;
      RECT 898.380 1.400 898.660 1617.000 ;
      RECT 900.620 1.400 900.900 1617.000 ;
      RECT 902.860 1.400 903.140 1617.000 ;
      RECT 905.100 1.400 905.380 1617.000 ;
      RECT 907.340 1.400 907.620 1617.000 ;
      RECT 909.580 1.400 909.860 1617.000 ;
      RECT 911.820 1.400 912.100 1617.000 ;
      RECT 914.060 1.400 914.340 1617.000 ;
      RECT 916.300 1.400 916.580 1617.000 ;
      RECT 918.540 1.400 918.820 1617.000 ;
      RECT 920.780 1.400 921.060 1617.000 ;
      RECT 923.020 1.400 923.300 1617.000 ;
      RECT 925.260 1.400 925.540 1617.000 ;
      RECT 927.500 1.400 927.780 1617.000 ;
      RECT 929.740 1.400 930.020 1617.000 ;
      RECT 931.980 1.400 932.260 1617.000 ;
      RECT 934.220 1.400 934.500 1617.000 ;
      RECT 936.460 1.400 936.740 1617.000 ;
      RECT 938.700 1.400 938.980 1617.000 ;
      RECT 940.940 1.400 941.220 1617.000 ;
      RECT 943.180 1.400 943.460 1617.000 ;
      RECT 945.420 1.400 945.700 1617.000 ;
      RECT 947.660 1.400 947.940 1617.000 ;
      RECT 949.900 1.400 950.180 1617.000 ;
      RECT 952.140 1.400 952.420 1617.000 ;
      RECT 954.380 1.400 954.660 1617.000 ;
      RECT 956.620 1.400 956.900 1617.000 ;
      RECT 958.860 1.400 959.140 1617.000 ;
      RECT 961.100 1.400 961.380 1617.000 ;
      RECT 963.340 1.400 963.620 1617.000 ;
      RECT 965.580 1.400 965.860 1617.000 ;
      RECT 967.820 1.400 968.100 1617.000 ;
      RECT 970.060 1.400 970.340 1617.000 ;
      RECT 972.300 1.400 972.580 1617.000 ;
      RECT 974.540 1.400 974.820 1617.000 ;
      RECT 976.780 1.400 977.060 1617.000 ;
      RECT 979.020 1.400 979.300 1617.000 ;
      RECT 981.260 1.400 981.540 1617.000 ;
      RECT 983.500 1.400 983.780 1617.000 ;
      RECT 985.740 1.400 986.020 1617.000 ;
      RECT 987.980 1.400 988.260 1617.000 ;
      RECT 990.220 1.400 990.500 1617.000 ;
      RECT 992.460 1.400 992.740 1617.000 ;
      RECT 994.700 1.400 994.980 1617.000 ;
      RECT 996.940 1.400 997.220 1617.000 ;
      RECT 999.180 1.400 999.460 1617.000 ;
      RECT 1001.420 1.400 1001.700 1617.000 ;
      RECT 1003.660 1.400 1003.940 1617.000 ;
      RECT 1005.900 1.400 1006.180 1617.000 ;
      RECT 1008.140 1.400 1008.420 1617.000 ;
      RECT 1010.380 1.400 1010.660 1617.000 ;
      RECT 1012.620 1.400 1012.900 1617.000 ;
      RECT 1014.860 1.400 1015.140 1617.000 ;
      RECT 1017.100 1.400 1017.380 1617.000 ;
      RECT 1019.340 1.400 1019.620 1617.000 ;
      RECT 1021.580 1.400 1021.860 1617.000 ;
      RECT 1023.820 1.400 1024.100 1617.000 ;
      RECT 1026.060 1.400 1026.340 1617.000 ;
      RECT 1028.300 1.400 1028.580 1617.000 ;
      RECT 1030.540 1.400 1030.820 1617.000 ;
      RECT 1032.780 1.400 1033.060 1617.000 ;
      RECT 1035.020 1.400 1035.300 1617.000 ;
      RECT 1037.260 1.400 1037.540 1617.000 ;
      RECT 1039.500 1.400 1039.780 1617.000 ;
      RECT 1041.740 1.400 1042.020 1617.000 ;
      RECT 1043.980 1.400 1044.260 1617.000 ;
      RECT 1046.220 1.400 1046.500 1617.000 ;
      RECT 1048.460 1.400 1048.740 1617.000 ;
      RECT 1050.700 1.400 1050.980 1617.000 ;
      RECT 1052.940 1.400 1053.220 1617.000 ;
      RECT 1055.180 1.400 1055.460 1617.000 ;
      RECT 1057.420 1.400 1057.700 1617.000 ;
      RECT 1059.660 1.400 1059.940 1617.000 ;
      RECT 1061.900 1.400 1062.180 1617.000 ;
      RECT 1064.140 1.400 1064.420 1617.000 ;
      RECT 1066.380 1.400 1066.660 1617.000 ;
      RECT 1068.620 1.400 1068.900 1617.000 ;
      RECT 1070.860 1.400 1071.140 1617.000 ;
      RECT 1073.100 1.400 1073.380 1617.000 ;
      RECT 1075.340 1.400 1075.620 1617.000 ;
      RECT 1077.580 1.400 1077.860 1617.000 ;
      RECT 1079.820 1.400 1080.100 1617.000 ;
      RECT 1082.060 1.400 1082.340 1617.000 ;
      RECT 1084.300 1.400 1084.580 1617.000 ;
      RECT 1086.540 1.400 1086.820 1617.000 ;
      RECT 1088.780 1.400 1089.060 1617.000 ;
      RECT 1091.020 1.400 1091.300 1617.000 ;
      RECT 1093.260 1.400 1093.540 1617.000 ;
      RECT 1095.500 1.400 1095.780 1617.000 ;
      RECT 1097.740 1.400 1098.020 1617.000 ;
      RECT 1099.980 1.400 1100.260 1617.000 ;
      RECT 1102.220 1.400 1102.500 1617.000 ;
      RECT 1104.460 1.400 1104.740 1617.000 ;
      RECT 1106.700 1.400 1106.980 1617.000 ;
      RECT 1108.940 1.400 1109.220 1617.000 ;
      RECT 1111.180 1.400 1111.460 1617.000 ;
      RECT 1113.420 1.400 1113.700 1617.000 ;
      RECT 1115.660 1.400 1115.940 1617.000 ;
      RECT 1117.900 1.400 1118.180 1617.000 ;
      RECT 1120.140 1.400 1120.420 1617.000 ;
      RECT 1122.380 1.400 1122.660 1617.000 ;
      RECT 1124.620 1.400 1124.900 1617.000 ;
      RECT 1126.860 1.400 1127.140 1617.000 ;
      RECT 1129.100 1.400 1129.380 1617.000 ;
      RECT 1131.340 1.400 1131.620 1617.000 ;
      RECT 1133.580 1.400 1133.860 1617.000 ;
      RECT 1135.820 1.400 1136.100 1617.000 ;
      RECT 1138.060 1.400 1138.340 1617.000 ;
      RECT 1140.300 1.400 1140.580 1617.000 ;
      RECT 1142.540 1.400 1142.820 1617.000 ;
      RECT 1144.780 1.400 1145.060 1617.000 ;
      RECT 1147.020 1.400 1147.300 1617.000 ;
      RECT 1149.260 1.400 1149.540 1617.000 ;
      RECT 1151.500 1.400 1151.780 1617.000 ;
      RECT 1153.740 1.400 1154.020 1617.000 ;
      RECT 1155.980 1.400 1156.260 1617.000 ;
      RECT 1158.220 1.400 1158.500 1617.000 ;
      RECT 1160.460 1.400 1160.740 1617.000 ;
      RECT 1162.700 1.400 1162.980 1617.000 ;
      RECT 1164.940 1.400 1165.220 1617.000 ;
      RECT 1167.180 1.400 1167.460 1617.000 ;
      RECT 1169.420 1.400 1169.700 1617.000 ;
      RECT 1171.660 1.400 1171.940 1617.000 ;
      RECT 1173.900 1.400 1174.180 1617.000 ;
      RECT 1176.140 1.400 1176.420 1617.000 ;
      RECT 1178.380 1.400 1178.660 1617.000 ;
      RECT 1180.620 1.400 1180.900 1617.000 ;
      RECT 1182.860 1.400 1183.140 1617.000 ;
      RECT 1185.100 1.400 1185.380 1617.000 ;
      RECT 1187.340 1.400 1187.620 1617.000 ;
      RECT 1189.580 1.400 1189.860 1617.000 ;
      RECT 1191.820 1.400 1192.100 1617.000 ;
      RECT 1194.060 1.400 1194.340 1617.000 ;
      RECT 1196.300 1.400 1196.580 1617.000 ;
      RECT 1198.540 1.400 1198.820 1617.000 ;
      RECT 1200.780 1.400 1201.060 1617.000 ;
      RECT 1203.020 1.400 1203.300 1617.000 ;
      RECT 1205.260 1.400 1205.540 1617.000 ;
      RECT 1207.500 1.400 1207.780 1617.000 ;
      RECT 1209.740 1.400 1210.020 1617.000 ;
      RECT 1211.980 1.400 1212.260 1617.000 ;
      RECT 1214.220 1.400 1214.500 1617.000 ;
      RECT 1216.460 1.400 1216.740 1617.000 ;
      RECT 1218.700 1.400 1218.980 1617.000 ;
      RECT 1220.940 1.400 1221.220 1617.000 ;
      RECT 1223.180 1.400 1223.460 1617.000 ;
      RECT 1225.420 1.400 1225.700 1617.000 ;
      RECT 1227.660 1.400 1227.940 1617.000 ;
      RECT 1229.900 1.400 1230.180 1617.000 ;
      RECT 1232.140 1.400 1232.420 1617.000 ;
      RECT 1234.380 1.400 1234.660 1617.000 ;
      RECT 1236.620 1.400 1236.900 1617.000 ;
      RECT 1238.860 1.400 1239.140 1617.000 ;
      RECT 1241.100 1.400 1241.380 1617.000 ;
      RECT 1243.340 1.400 1243.620 1617.000 ;
      RECT 1245.580 1.400 1245.860 1617.000 ;
      RECT 1247.820 1.400 1248.100 1617.000 ;
      RECT 1250.060 1.400 1250.340 1617.000 ;
      RECT 1252.300 1.400 1252.580 1617.000 ;
      RECT 1254.540 1.400 1254.820 1617.000 ;
      RECT 1256.780 1.400 1257.060 1617.000 ;
      RECT 1259.020 1.400 1259.300 1617.000 ;
      RECT 1261.260 1.400 1261.540 1617.000 ;
      RECT 1263.500 1.400 1263.780 1617.000 ;
      RECT 1265.740 1.400 1266.020 1617.000 ;
      RECT 1267.980 1.400 1268.260 1617.000 ;
      RECT 1270.220 1.400 1270.500 1617.000 ;
      RECT 1272.460 1.400 1272.740 1617.000 ;
      RECT 1274.700 1.400 1274.980 1617.000 ;
      RECT 1276.940 1.400 1277.220 1617.000 ;
      RECT 1279.180 1.400 1279.460 1617.000 ;
      RECT 1281.420 1.400 1281.700 1617.000 ;
      RECT 1283.660 1.400 1283.940 1617.000 ;
      RECT 1285.900 1.400 1286.180 1617.000 ;
      RECT 1288.140 1.400 1288.420 1617.000 ;
      RECT 1290.380 1.400 1290.660 1617.000 ;
      RECT 1292.620 1.400 1292.900 1617.000 ;
      RECT 1294.860 1.400 1295.140 1617.000 ;
      RECT 1297.100 1.400 1297.380 1617.000 ;
      RECT 1299.340 1.400 1299.620 1617.000 ;
      RECT 1301.580 1.400 1301.860 1617.000 ;
      RECT 1303.820 1.400 1304.100 1617.000 ;
      RECT 1306.060 1.400 1306.340 1617.000 ;
      RECT 1308.300 1.400 1308.580 1617.000 ;
      RECT 1310.540 1.400 1310.820 1617.000 ;
      RECT 1312.780 1.400 1313.060 1617.000 ;
      RECT 1315.020 1.400 1315.300 1617.000 ;
      RECT 1317.260 1.400 1317.540 1617.000 ;
      RECT 1319.500 1.400 1319.780 1617.000 ;
      RECT 1321.740 1.400 1322.020 1617.000 ;
      RECT 1323.980 1.400 1324.260 1617.000 ;
      RECT 1326.220 1.400 1326.500 1617.000 ;
      RECT 1328.460 1.400 1328.740 1617.000 ;
      RECT 1330.700 1.400 1330.980 1617.000 ;
      RECT 1332.940 1.400 1333.220 1617.000 ;
      RECT 1335.180 1.400 1335.460 1617.000 ;
      RECT 1337.420 1.400 1337.700 1617.000 ;
      RECT 1339.660 1.400 1339.940 1617.000 ;
      RECT 1341.900 1.400 1342.180 1617.000 ;
      RECT 1344.140 1.400 1344.420 1617.000 ;
      RECT 1346.380 1.400 1346.660 1617.000 ;
      RECT 1348.620 1.400 1348.900 1617.000 ;
      RECT 1350.860 1.400 1351.140 1617.000 ;
      RECT 1353.100 1.400 1353.380 1617.000 ;
      RECT 1355.340 1.400 1355.620 1617.000 ;
      RECT 1357.580 1.400 1357.860 1617.000 ;
      RECT 1359.820 1.400 1360.100 1617.000 ;
      RECT 1362.060 1.400 1362.340 1617.000 ;
      RECT 1364.300 1.400 1364.580 1617.000 ;
      RECT 1366.540 1.400 1366.820 1617.000 ;
      RECT 1368.780 1.400 1369.060 1617.000 ;
      RECT 1371.020 1.400 1371.300 1617.000 ;
      RECT 1373.260 1.400 1373.540 1617.000 ;
      RECT 1375.500 1.400 1375.780 1617.000 ;
      RECT 1377.740 1.400 1378.020 1617.000 ;
      RECT 1379.980 1.400 1380.260 1617.000 ;
      RECT 1382.220 1.400 1382.500 1617.000 ;
      RECT 1384.460 1.400 1384.740 1617.000 ;
      RECT 1386.700 1.400 1386.980 1617.000 ;
      RECT 1388.940 1.400 1389.220 1617.000 ;
      RECT 1391.180 1.400 1391.460 1617.000 ;
      RECT 1393.420 1.400 1393.700 1617.000 ;
      RECT 1395.660 1.400 1395.940 1617.000 ;
      RECT 1397.900 1.400 1398.180 1617.000 ;
      RECT 1400.140 1.400 1400.420 1617.000 ;
      RECT 1402.380 1.400 1402.660 1617.000 ;
      RECT 1404.620 1.400 1404.900 1617.000 ;
      RECT 1406.860 1.400 1407.140 1617.000 ;
      RECT 1409.100 1.400 1409.380 1617.000 ;
      RECT 1411.340 1.400 1411.620 1617.000 ;
      RECT 1413.580 1.400 1413.860 1617.000 ;
      RECT 1415.820 1.400 1416.100 1617.000 ;
      RECT 1418.060 1.400 1418.340 1617.000 ;
      RECT 1420.300 1.400 1420.580 1617.000 ;
      RECT 1422.540 1.400 1422.820 1617.000 ;
      RECT 1424.780 1.400 1425.060 1617.000 ;
      RECT 1427.020 1.400 1427.300 1617.000 ;
      RECT 1429.260 1.400 1429.540 1617.000 ;
      RECT 1431.500 1.400 1431.780 1617.000 ;
      RECT 1433.740 1.400 1434.020 1617.000 ;
      RECT 1435.980 1.400 1436.260 1617.000 ;
      RECT 1438.220 1.400 1438.500 1617.000 ;
      RECT 1440.460 1.400 1440.740 1617.000 ;
      RECT 1442.700 1.400 1442.980 1617.000 ;
      RECT 1444.940 1.400 1445.220 1617.000 ;
      RECT 1447.180 1.400 1447.460 1617.000 ;
      RECT 1449.420 1.400 1449.700 1617.000 ;
      RECT 1451.660 1.400 1451.940 1617.000 ;
      RECT 1453.900 1.400 1454.180 1617.000 ;
      RECT 1456.140 1.400 1456.420 1617.000 ;
      RECT 1458.380 1.400 1458.660 1617.000 ;
      RECT 1460.620 1.400 1460.900 1617.000 ;
      RECT 1462.860 1.400 1463.140 1617.000 ;
      RECT 1465.100 1.400 1465.380 1617.000 ;
      RECT 1467.340 1.400 1467.620 1617.000 ;
      RECT 1469.580 1.400 1469.860 1617.000 ;
      RECT 1471.820 1.400 1472.100 1617.000 ;
      RECT 1474.060 1.400 1474.340 1617.000 ;
      RECT 1476.300 1.400 1476.580 1617.000 ;
      RECT 1478.540 1.400 1478.820 1617.000 ;
      RECT 1480.780 1.400 1481.060 1617.000 ;
      RECT 1483.020 1.400 1483.300 1617.000 ;
      RECT 1485.260 1.400 1485.540 1617.000 ;
      RECT 1487.500 1.400 1487.780 1617.000 ;
      RECT 1489.740 1.400 1490.020 1617.000 ;
      RECT 1491.980 1.400 1492.260 1617.000 ;
      RECT 1494.220 1.400 1494.500 1617.000 ;
      RECT 1496.460 1.400 1496.740 1617.000 ;
      RECT 1498.700 1.400 1498.980 1617.000 ;
      RECT 1500.940 1.400 1501.220 1617.000 ;
      RECT 1503.180 1.400 1503.460 1617.000 ;
      RECT 1505.420 1.400 1505.700 1617.000 ;
      RECT 1507.660 1.400 1507.940 1617.000 ;
      RECT 1509.900 1.400 1510.180 1617.000 ;
      RECT 1512.140 1.400 1512.420 1617.000 ;
      RECT 1514.380 1.400 1514.660 1617.000 ;
      RECT 1516.620 1.400 1516.900 1617.000 ;
      RECT 1518.860 1.400 1519.140 1617.000 ;
      RECT 1521.100 1.400 1521.380 1617.000 ;
      RECT 1523.340 1.400 1523.620 1617.000 ;
      RECT 1525.580 1.400 1525.860 1617.000 ;
      RECT 1527.820 1.400 1528.100 1617.000 ;
      RECT 1530.060 1.400 1530.340 1617.000 ;
      RECT 1532.300 1.400 1532.580 1617.000 ;
      RECT 1534.540 1.400 1534.820 1617.000 ;
      RECT 1536.780 1.400 1537.060 1617.000 ;
      RECT 1539.020 1.400 1539.300 1617.000 ;
      RECT 1541.260 1.400 1541.540 1617.000 ;
      RECT 1543.500 1.400 1543.780 1617.000 ;
      RECT 1545.740 1.400 1546.020 1617.000 ;
      RECT 1547.980 1.400 1548.260 1617.000 ;
      RECT 1550.220 1.400 1550.500 1617.000 ;
      RECT 1552.460 1.400 1552.740 1617.000 ;
      RECT 1554.700 1.400 1554.980 1617.000 ;
      RECT 1556.940 1.400 1557.220 1617.000 ;
      RECT 1559.180 1.400 1559.460 1617.000 ;
      RECT 1561.420 1.400 1561.700 1617.000 ;
      RECT 1563.660 1.400 1563.940 1617.000 ;
      RECT 1565.900 1.400 1566.180 1617.000 ;
      RECT 1568.140 1.400 1568.420 1617.000 ;
      RECT 1570.380 1.400 1570.660 1617.000 ;
      RECT 1572.620 1.400 1572.900 1617.000 ;
      RECT 1574.860 1.400 1575.140 1617.000 ;
      RECT 1577.100 1.400 1577.380 1617.000 ;
      RECT 1579.340 1.400 1579.620 1617.000 ;
      RECT 1581.580 1.400 1581.860 1617.000 ;
      RECT 1583.820 1.400 1584.100 1617.000 ;
      RECT 1586.060 1.400 1586.340 1617.000 ;
      RECT 1588.300 1.400 1588.580 1617.000 ;
      RECT 1590.540 1.400 1590.820 1617.000 ;
      RECT 1592.780 1.400 1593.060 1617.000 ;
      RECT 1595.020 1.400 1595.300 1617.000 ;
      RECT 1597.260 1.400 1597.540 1617.000 ;
      RECT 1599.500 1.400 1599.780 1617.000 ;
      RECT 1601.740 1.400 1602.020 1617.000 ;
      RECT 1603.980 1.400 1604.260 1617.000 ;
      RECT 1606.220 1.400 1606.500 1617.000 ;
      RECT 1608.460 1.400 1608.740 1617.000 ;
      RECT 1610.700 1.400 1610.980 1617.000 ;
      RECT 1612.940 1.400 1613.220 1617.000 ;
      RECT 1615.180 1.400 1615.460 1617.000 ;
      RECT 1617.420 1.400 1617.700 1617.000 ;
      RECT 1619.660 1.400 1619.940 1617.000 ;
      RECT 1621.900 1.400 1622.180 1617.000 ;
      RECT 1624.140 1.400 1624.420 1617.000 ;
      RECT 1626.380 1.400 1626.660 1617.000 ;
      RECT 1628.620 1.400 1628.900 1617.000 ;
      RECT 1630.860 1.400 1631.140 1617.000 ;
      RECT 1633.100 1.400 1633.380 1617.000 ;
      RECT 1635.340 1.400 1635.620 1617.000 ;
      RECT 1637.580 1.400 1637.860 1617.000 ;
      RECT 1639.820 1.400 1640.100 1617.000 ;
      RECT 1642.060 1.400 1642.340 1617.000 ;
      RECT 1644.300 1.400 1644.580 1617.000 ;
      RECT 1646.540 1.400 1646.820 1617.000 ;
      RECT 1648.780 1.400 1649.060 1617.000 ;
      RECT 1651.020 1.400 1651.300 1617.000 ;
      RECT 1653.260 1.400 1653.540 1617.000 ;
      RECT 1655.500 1.400 1655.780 1617.000 ;
      RECT 1657.740 1.400 1658.020 1617.000 ;
      RECT 1659.980 1.400 1660.260 1617.000 ;
      RECT 1662.220 1.400 1662.500 1617.000 ;
      RECT 1664.460 1.400 1664.740 1617.000 ;
      RECT 1666.700 1.400 1666.980 1617.000 ;
      RECT 1668.940 1.400 1669.220 1617.000 ;
      RECT 1671.180 1.400 1671.460 1617.000 ;
      RECT 1673.420 1.400 1673.700 1617.000 ;
      RECT 1675.660 1.400 1675.940 1617.000 ;
      RECT 1677.900 1.400 1678.180 1617.000 ;
      RECT 1680.140 1.400 1680.420 1617.000 ;
      RECT 1682.380 1.400 1682.660 1617.000 ;
      RECT 1684.620 1.400 1684.900 1617.000 ;
      RECT 1686.860 1.400 1687.140 1617.000 ;
      RECT 1689.100 1.400 1689.380 1617.000 ;
      RECT 1691.340 1.400 1691.620 1617.000 ;
      RECT 1693.580 1.400 1693.860 1617.000 ;
      RECT 1695.820 1.400 1696.100 1617.000 ;
      RECT 1698.060 1.400 1698.340 1617.000 ;
      RECT 1700.300 1.400 1700.580 1617.000 ;
      RECT 1702.540 1.400 1702.820 1617.000 ;
      RECT 1704.780 1.400 1705.060 1617.000 ;
      RECT 1707.020 1.400 1707.300 1617.000 ;
      RECT 1709.260 1.400 1709.540 1617.000 ;
      RECT 1711.500 1.400 1711.780 1617.000 ;
      RECT 1713.740 1.400 1714.020 1617.000 ;
      RECT 1715.980 1.400 1716.260 1617.000 ;
      RECT 1718.220 1.400 1718.500 1617.000 ;
      RECT 1720.460 1.400 1720.740 1617.000 ;
      RECT 1722.700 1.400 1722.980 1617.000 ;
      RECT 1724.940 1.400 1725.220 1617.000 ;
      RECT 1727.180 1.400 1727.460 1617.000 ;
      RECT 1729.420 1.400 1729.700 1617.000 ;
      RECT 1731.660 1.400 1731.940 1617.000 ;
      RECT 1733.900 1.400 1734.180 1617.000 ;
      RECT 1736.140 1.400 1736.420 1617.000 ;
      RECT 1738.380 1.400 1738.660 1617.000 ;
      RECT 1740.620 1.400 1740.900 1617.000 ;
      RECT 1742.860 1.400 1743.140 1617.000 ;
      RECT 1745.100 1.400 1745.380 1617.000 ;
      RECT 1747.340 1.400 1747.620 1617.000 ;
      RECT 1749.580 1.400 1749.860 1617.000 ;
      RECT 1751.820 1.400 1752.100 1617.000 ;
      RECT 1754.060 1.400 1754.340 1617.000 ;
      RECT 1756.300 1.400 1756.580 1617.000 ;
      RECT 1758.540 1.400 1758.820 1617.000 ;
      RECT 1760.780 1.400 1761.060 1617.000 ;
      RECT 1763.020 1.400 1763.300 1617.000 ;
      RECT 1765.260 1.400 1765.540 1617.000 ;
      RECT 1767.500 1.400 1767.780 1617.000 ;
      RECT 1769.740 1.400 1770.020 1617.000 ;
      RECT 1771.980 1.400 1772.260 1617.000 ;
      RECT 1774.220 1.400 1774.500 1617.000 ;
      RECT 1776.460 1.400 1776.740 1617.000 ;
      RECT 1778.700 1.400 1778.980 1617.000 ;
      RECT 1780.940 1.400 1781.220 1617.000 ;
      RECT 1783.180 1.400 1783.460 1617.000 ;
      RECT 1785.420 1.400 1785.700 1617.000 ;
      RECT 1787.660 1.400 1787.940 1617.000 ;
      RECT 1789.900 1.400 1790.180 1617.000 ;
      RECT 1792.140 1.400 1792.420 1617.000 ;
      RECT 1794.380 1.400 1794.660 1617.000 ;
      RECT 1796.620 1.400 1796.900 1617.000 ;
      RECT 1798.860 1.400 1799.140 1617.000 ;
      RECT 1801.100 1.400 1801.380 1617.000 ;
      RECT 1803.340 1.400 1803.620 1617.000 ;
      RECT 1805.580 1.400 1805.860 1617.000 ;
      RECT 1807.820 1.400 1808.100 1617.000 ;
      RECT 1810.060 1.400 1810.340 1617.000 ;
      RECT 1812.300 1.400 1812.580 1617.000 ;
      RECT 1814.540 1.400 1814.820 1617.000 ;
      RECT 1816.780 1.400 1817.060 1617.000 ;
      RECT 1819.020 1.400 1819.300 1617.000 ;
      RECT 1821.260 1.400 1821.540 1617.000 ;
      RECT 1823.500 1.400 1823.780 1617.000 ;
      RECT 1825.740 1.400 1826.020 1617.000 ;
      RECT 1827.980 1.400 1828.260 1617.000 ;
      RECT 1830.220 1.400 1830.500 1617.000 ;
      RECT 1832.460 1.400 1832.740 1617.000 ;
      RECT 1834.700 1.400 1834.980 1617.000 ;
      RECT 1836.940 1.400 1837.220 1617.000 ;
      RECT 1839.180 1.400 1839.460 1617.000 ;
      RECT 1841.420 1.400 1841.700 1617.000 ;
      RECT 1843.660 1.400 1843.940 1617.000 ;
      RECT 1845.900 1.400 1846.180 1617.000 ;
      RECT 1848.140 1.400 1848.420 1617.000 ;
      RECT 1850.380 1.400 1850.660 1617.000 ;
      RECT 1852.620 1.400 1852.900 1617.000 ;
      RECT 1854.860 1.400 1855.140 1617.000 ;
      RECT 1857.100 1.400 1857.380 1617.000 ;
      RECT 1859.340 1.400 1859.620 1617.000 ;
      RECT 1861.580 1.400 1861.860 1617.000 ;
      RECT 1863.820 1.400 1864.100 1617.000 ;
      RECT 1866.060 1.400 1866.340 1617.000 ;
      RECT 1868.300 1.400 1868.580 1617.000 ;
      RECT 1870.540 1.400 1870.820 1617.000 ;
      RECT 1872.780 1.400 1873.060 1617.000 ;
      RECT 1875.020 1.400 1875.300 1617.000 ;
      RECT 1877.260 1.400 1877.540 1617.000 ;
      RECT 1879.500 1.400 1879.780 1617.000 ;
      RECT 1881.740 1.400 1882.020 1617.000 ;
      RECT 1883.980 1.400 1884.260 1617.000 ;
      RECT 1886.220 1.400 1886.500 1617.000 ;
      RECT 1888.460 1.400 1888.740 1617.000 ;
      RECT 1890.700 1.400 1890.980 1617.000 ;
      RECT 1892.940 1.400 1893.220 1617.000 ;
      RECT 1895.180 1.400 1895.460 1617.000 ;
      RECT 1897.420 1.400 1897.700 1617.000 ;
      RECT 1899.660 1.400 1899.940 1617.000 ;
      RECT 1901.900 1.400 1902.180 1617.000 ;
      RECT 1904.140 1.400 1904.420 1617.000 ;
      RECT 1906.380 1.400 1906.660 1617.000 ;
      RECT 1908.620 1.400 1908.900 1617.000 ;
      RECT 1910.860 1.400 1911.140 1617.000 ;
      RECT 1913.100 1.400 1913.380 1617.000 ;
      RECT 1915.340 1.400 1915.620 1617.000 ;
      RECT 1917.580 1.400 1917.860 1617.000 ;
      RECT 1919.820 1.400 1920.100 1617.000 ;
      RECT 1922.060 1.400 1922.340 1617.000 ;
      RECT 1924.300 1.400 1924.580 1617.000 ;
      RECT 1926.540 1.400 1926.820 1617.000 ;
      RECT 1928.780 1.400 1929.060 1617.000 ;
      RECT 1931.020 1.400 1931.300 1617.000 ;
      RECT 1933.260 1.400 1933.540 1617.000 ;
      RECT 1935.500 1.400 1935.780 1617.000 ;
      RECT 1937.740 1.400 1938.020 1617.000 ;
      RECT 1939.980 1.400 1940.260 1617.000 ;
      RECT 1942.220 1.400 1942.500 1617.000 ;
      RECT 1944.460 1.400 1944.740 1617.000 ;
      RECT 1946.700 1.400 1946.980 1617.000 ;
      RECT 1948.940 1.400 1949.220 1617.000 ;
      RECT 1951.180 1.400 1951.460 1617.000 ;
      RECT 1953.420 1.400 1953.700 1617.000 ;
      RECT 1955.660 1.400 1955.940 1617.000 ;
      RECT 1957.900 1.400 1958.180 1617.000 ;
      RECT 1960.140 1.400 1960.420 1617.000 ;
      RECT 1962.380 1.400 1962.660 1617.000 ;
      RECT 1964.620 1.400 1964.900 1617.000 ;
      RECT 1966.860 1.400 1967.140 1617.000 ;
      RECT 1969.100 1.400 1969.380 1617.000 ;
      RECT 1971.340 1.400 1971.620 1617.000 ;
      RECT 1973.580 1.400 1973.860 1617.000 ;
      RECT 1975.820 1.400 1976.100 1617.000 ;
      RECT 1978.060 1.400 1978.340 1617.000 ;
      RECT 1980.300 1.400 1980.580 1617.000 ;
      RECT 1982.540 1.400 1982.820 1617.000 ;
      RECT 1984.780 1.400 1985.060 1617.000 ;
      RECT 1987.020 1.400 1987.300 1617.000 ;
      RECT 1989.260 1.400 1989.540 1617.000 ;
      RECT 1991.500 1.400 1991.780 1617.000 ;
      RECT 1993.740 1.400 1994.020 1617.000 ;
      RECT 1995.980 1.400 1996.260 1617.000 ;
      RECT 1998.220 1.400 1998.500 1617.000 ;
      RECT 2000.460 1.400 2000.740 1617.000 ;
      RECT 2002.700 1.400 2002.980 1617.000 ;
      RECT 2004.940 1.400 2005.220 1617.000 ;
      RECT 2007.180 1.400 2007.460 1617.000 ;
      RECT 2009.420 1.400 2009.700 1617.000 ;
      RECT 2011.660 1.400 2011.940 1617.000 ;
      RECT 2013.900 1.400 2014.180 1617.000 ;
      RECT 2016.140 1.400 2016.420 1617.000 ;
      RECT 2018.380 1.400 2018.660 1617.000 ;
      RECT 2020.620 1.400 2020.900 1617.000 ;
      RECT 2022.860 1.400 2023.140 1617.000 ;
      RECT 2025.100 1.400 2025.380 1617.000 ;
      RECT 2027.340 1.400 2027.620 1617.000 ;
      RECT 2029.580 1.400 2029.860 1617.000 ;
      RECT 2031.820 1.400 2032.100 1617.000 ;
      RECT 2034.060 1.400 2034.340 1617.000 ;
      RECT 2036.300 1.400 2036.580 1617.000 ;
      RECT 2038.540 1.400 2038.820 1617.000 ;
      RECT 2040.780 1.400 2041.060 1617.000 ;
      RECT 2043.020 1.400 2043.300 1617.000 ;
      RECT 2045.260 1.400 2045.540 1617.000 ;
      RECT 2047.500 1.400 2047.780 1617.000 ;
      RECT 2049.740 1.400 2050.020 1617.000 ;
      RECT 2051.980 1.400 2052.260 1617.000 ;
      RECT 2054.220 1.400 2054.500 1617.000 ;
      RECT 2056.460 1.400 2056.740 1617.000 ;
      RECT 2058.700 1.400 2058.980 1617.000 ;
      RECT 2060.940 1.400 2061.220 1617.000 ;
      RECT 2063.180 1.400 2063.460 1617.000 ;
      RECT 2065.420 1.400 2065.700 1617.000 ;
      RECT 2067.660 1.400 2067.940 1617.000 ;
      RECT 2069.900 1.400 2070.180 1617.000 ;
      RECT 2072.140 1.400 2072.420 1617.000 ;
      RECT 2074.380 1.400 2074.660 1617.000 ;
      RECT 2076.620 1.400 2076.900 1617.000 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 2078.600 1618.400 ;
    LAYER metal2 ;
    RECT 0 0 2078.600 1618.400 ;
    LAYER metal3 ;
    RECT 0.070 0 2078.600 1618.400 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.505 ;
    RECT 0 1.575 0.070 1.645 ;
    RECT 0 1.715 0.070 1.785 ;
    RECT 0 1.855 0.070 1.925 ;
    RECT 0 1.995 0.070 2.065 ;
    RECT 0 2.135 0.070 2.205 ;
    RECT 0 2.275 0.070 2.345 ;
    RECT 0 2.415 0.070 2.485 ;
    RECT 0 2.555 0.070 2.625 ;
    RECT 0 2.695 0.070 2.765 ;
    RECT 0 2.835 0.070 2.905 ;
    RECT 0 2.975 0.070 3.045 ;
    RECT 0 3.115 0.070 3.185 ;
    RECT 0 3.255 0.070 3.325 ;
    RECT 0 3.395 0.070 3.465 ;
    RECT 0 3.535 0.070 3.605 ;
    RECT 0 3.675 0.070 3.745 ;
    RECT 0 3.815 0.070 3.885 ;
    RECT 0 3.955 0.070 4.025 ;
    RECT 0 4.095 0.070 4.165 ;
    RECT 0 4.235 0.070 4.305 ;
    RECT 0 4.375 0.070 4.445 ;
    RECT 0 4.515 0.070 4.585 ;
    RECT 0 4.655 0.070 4.725 ;
    RECT 0 4.795 0.070 4.865 ;
    RECT 0 4.935 0.070 5.005 ;
    RECT 0 5.075 0.070 5.145 ;
    RECT 0 5.215 0.070 5.285 ;
    RECT 0 5.355 0.070 5.425 ;
    RECT 0 5.495 0.070 5.565 ;
    RECT 0 5.635 0.070 5.705 ;
    RECT 0 5.775 0.070 5.845 ;
    RECT 0 5.915 0.070 5.985 ;
    RECT 0 6.055 0.070 6.125 ;
    RECT 0 6.195 0.070 6.265 ;
    RECT 0 6.335 0.070 6.405 ;
    RECT 0 6.475 0.070 6.545 ;
    RECT 0 6.615 0.070 6.685 ;
    RECT 0 6.755 0.070 6.825 ;
    RECT 0 6.895 0.070 6.965 ;
    RECT 0 7.035 0.070 7.105 ;
    RECT 0 7.175 0.070 7.245 ;
    RECT 0 7.315 0.070 7.385 ;
    RECT 0 7.455 0.070 7.525 ;
    RECT 0 7.595 0.070 7.665 ;
    RECT 0 7.735 0.070 7.805 ;
    RECT 0 7.875 0.070 7.945 ;
    RECT 0 8.015 0.070 8.085 ;
    RECT 0 8.155 0.070 8.225 ;
    RECT 0 8.295 0.070 8.365 ;
    RECT 0 8.435 0.070 8.505 ;
    RECT 0 8.575 0.070 8.645 ;
    RECT 0 8.715 0.070 8.785 ;
    RECT 0 8.855 0.070 8.925 ;
    RECT 0 8.995 0.070 9.065 ;
    RECT 0 9.135 0.070 9.205 ;
    RECT 0 9.275 0.070 9.345 ;
    RECT 0 9.415 0.070 9.485 ;
    RECT 0 9.555 0.070 9.625 ;
    RECT 0 9.695 0.070 9.765 ;
    RECT 0 9.835 0.070 9.905 ;
    RECT 0 9.975 0.070 10.045 ;
    RECT 0 10.115 0.070 10.185 ;
    RECT 0 10.255 0.070 10.325 ;
    RECT 0 10.395 0.070 10.465 ;
    RECT 0 10.535 0.070 10.605 ;
    RECT 0 10.675 0.070 10.745 ;
    RECT 0 10.815 0.070 10.885 ;
    RECT 0 10.955 0.070 11.025 ;
    RECT 0 11.095 0.070 11.165 ;
    RECT 0 11.235 0.070 11.305 ;
    RECT 0 11.375 0.070 11.445 ;
    RECT 0 11.515 0.070 11.585 ;
    RECT 0 11.655 0.070 11.725 ;
    RECT 0 11.795 0.070 11.865 ;
    RECT 0 11.935 0.070 12.005 ;
    RECT 0 12.075 0.070 12.145 ;
    RECT 0 12.215 0.070 12.285 ;
    RECT 0 12.355 0.070 12.425 ;
    RECT 0 12.495 0.070 12.565 ;
    RECT 0 12.635 0.070 12.705 ;
    RECT 0 12.775 0.070 12.845 ;
    RECT 0 12.915 0.070 12.985 ;
    RECT 0 13.055 0.070 13.125 ;
    RECT 0 13.195 0.070 13.265 ;
    RECT 0 13.335 0.070 13.405 ;
    RECT 0 13.475 0.070 13.545 ;
    RECT 0 13.615 0.070 13.685 ;
    RECT 0 13.755 0.070 13.825 ;
    RECT 0 13.895 0.070 13.965 ;
    RECT 0 14.035 0.070 14.105 ;
    RECT 0 14.175 0.070 14.245 ;
    RECT 0 14.315 0.070 14.385 ;
    RECT 0 14.455 0.070 14.525 ;
    RECT 0 14.595 0.070 14.665 ;
    RECT 0 14.735 0.070 14.805 ;
    RECT 0 14.875 0.070 14.945 ;
    RECT 0 15.015 0.070 15.085 ;
    RECT 0 15.155 0.070 15.225 ;
    RECT 0 15.295 0.070 15.365 ;
    RECT 0 15.435 0.070 15.505 ;
    RECT 0 15.575 0.070 15.645 ;
    RECT 0 15.715 0.070 15.785 ;
    RECT 0 15.855 0.070 15.925 ;
    RECT 0 15.995 0.070 16.065 ;
    RECT 0 16.135 0.070 16.205 ;
    RECT 0 16.275 0.070 16.345 ;
    RECT 0 16.415 0.070 16.485 ;
    RECT 0 16.555 0.070 16.625 ;
    RECT 0 16.695 0.070 16.765 ;
    RECT 0 16.835 0.070 16.905 ;
    RECT 0 16.975 0.070 17.045 ;
    RECT 0 17.115 0.070 17.185 ;
    RECT 0 17.255 0.070 17.325 ;
    RECT 0 17.395 0.070 17.465 ;
    RECT 0 17.535 0.070 17.605 ;
    RECT 0 17.675 0.070 17.745 ;
    RECT 0 17.815 0.070 17.885 ;
    RECT 0 17.955 0.070 18.025 ;
    RECT 0 18.095 0.070 18.165 ;
    RECT 0 18.235 0.070 18.305 ;
    RECT 0 18.375 0.070 18.445 ;
    RECT 0 18.515 0.070 18.585 ;
    RECT 0 18.655 0.070 18.725 ;
    RECT 0 18.795 0.070 18.865 ;
    RECT 0 18.935 0.070 19.005 ;
    RECT 0 19.075 0.070 19.145 ;
    RECT 0 19.215 0.070 19.285 ;
    RECT 0 19.355 0.070 19.425 ;
    RECT 0 19.495 0.070 19.565 ;
    RECT 0 19.635 0.070 19.705 ;
    RECT 0 19.775 0.070 19.845 ;
    RECT 0 19.915 0.070 19.985 ;
    RECT 0 20.055 0.070 20.125 ;
    RECT 0 20.195 0.070 20.265 ;
    RECT 0 20.335 0.070 20.405 ;
    RECT 0 20.475 0.070 20.545 ;
    RECT 0 20.615 0.070 20.685 ;
    RECT 0 20.755 0.070 20.825 ;
    RECT 0 20.895 0.070 20.965 ;
    RECT 0 21.035 0.070 21.105 ;
    RECT 0 21.175 0.070 21.245 ;
    RECT 0 21.315 0.070 21.385 ;
    RECT 0 21.455 0.070 21.525 ;
    RECT 0 21.595 0.070 21.665 ;
    RECT 0 21.735 0.070 21.805 ;
    RECT 0 21.875 0.070 21.945 ;
    RECT 0 22.015 0.070 22.085 ;
    RECT 0 22.155 0.070 22.225 ;
    RECT 0 22.295 0.070 22.365 ;
    RECT 0 22.435 0.070 22.505 ;
    RECT 0 22.575 0.070 22.645 ;
    RECT 0 22.715 0.070 22.785 ;
    RECT 0 22.855 0.070 22.925 ;
    RECT 0 22.995 0.070 23.065 ;
    RECT 0 23.135 0.070 23.205 ;
    RECT 0 23.275 0.070 23.345 ;
    RECT 0 23.415 0.070 23.485 ;
    RECT 0 23.555 0.070 23.625 ;
    RECT 0 23.695 0.070 23.765 ;
    RECT 0 23.835 0.070 23.905 ;
    RECT 0 23.975 0.070 24.045 ;
    RECT 0 24.115 0.070 24.185 ;
    RECT 0 24.255 0.070 24.325 ;
    RECT 0 24.395 0.070 24.465 ;
    RECT 0 24.535 0.070 24.605 ;
    RECT 0 24.675 0.070 24.745 ;
    RECT 0 24.815 0.070 24.885 ;
    RECT 0 24.955 0.070 25.025 ;
    RECT 0 25.095 0.070 25.165 ;
    RECT 0 25.235 0.070 25.305 ;
    RECT 0 25.375 0.070 25.445 ;
    RECT 0 25.515 0.070 25.585 ;
    RECT 0 25.655 0.070 25.725 ;
    RECT 0 25.795 0.070 25.865 ;
    RECT 0 25.935 0.070 26.005 ;
    RECT 0 26.075 0.070 26.145 ;
    RECT 0 26.215 0.070 26.285 ;
    RECT 0 26.355 0.070 26.425 ;
    RECT 0 26.495 0.070 26.565 ;
    RECT 0 26.635 0.070 26.705 ;
    RECT 0 26.775 0.070 26.845 ;
    RECT 0 26.915 0.070 26.985 ;
    RECT 0 27.055 0.070 27.125 ;
    RECT 0 27.195 0.070 27.265 ;
    RECT 0 27.335 0.070 27.405 ;
    RECT 0 27.475 0.070 27.545 ;
    RECT 0 27.615 0.070 27.685 ;
    RECT 0 27.755 0.070 27.825 ;
    RECT 0 27.895 0.070 27.965 ;
    RECT 0 28.035 0.070 28.105 ;
    RECT 0 28.175 0.070 28.245 ;
    RECT 0 28.315 0.070 28.385 ;
    RECT 0 28.455 0.070 28.525 ;
    RECT 0 28.595 0.070 28.665 ;
    RECT 0 28.735 0.070 28.805 ;
    RECT 0 28.875 0.070 28.945 ;
    RECT 0 29.015 0.070 29.085 ;
    RECT 0 29.155 0.070 29.225 ;
    RECT 0 29.295 0.070 29.365 ;
    RECT 0 29.435 0.070 29.505 ;
    RECT 0 29.575 0.070 29.645 ;
    RECT 0 29.715 0.070 29.785 ;
    RECT 0 29.855 0.070 29.925 ;
    RECT 0 29.995 0.070 30.065 ;
    RECT 0 30.135 0.070 30.205 ;
    RECT 0 30.275 0.070 30.345 ;
    RECT 0 30.415 0.070 30.485 ;
    RECT 0 30.555 0.070 30.625 ;
    RECT 0 30.695 0.070 30.765 ;
    RECT 0 30.835 0.070 30.905 ;
    RECT 0 30.975 0.070 31.045 ;
    RECT 0 31.115 0.070 31.185 ;
    RECT 0 31.255 0.070 31.325 ;
    RECT 0 31.395 0.070 31.465 ;
    RECT 0 31.535 0.070 31.605 ;
    RECT 0 31.675 0.070 31.745 ;
    RECT 0 31.815 0.070 31.885 ;
    RECT 0 31.955 0.070 32.025 ;
    RECT 0 32.095 0.070 32.165 ;
    RECT 0 32.235 0.070 32.305 ;
    RECT 0 32.375 0.070 32.445 ;
    RECT 0 32.515 0.070 32.585 ;
    RECT 0 32.655 0.070 32.725 ;
    RECT 0 32.795 0.070 32.865 ;
    RECT 0 32.935 0.070 33.005 ;
    RECT 0 33.075 0.070 33.145 ;
    RECT 0 33.215 0.070 33.285 ;
    RECT 0 33.355 0.070 33.425 ;
    RECT 0 33.495 0.070 33.565 ;
    RECT 0 33.635 0.070 33.705 ;
    RECT 0 33.775 0.070 33.845 ;
    RECT 0 33.915 0.070 33.985 ;
    RECT 0 34.055 0.070 34.125 ;
    RECT 0 34.195 0.070 34.265 ;
    RECT 0 34.335 0.070 34.405 ;
    RECT 0 34.475 0.070 34.545 ;
    RECT 0 34.615 0.070 34.685 ;
    RECT 0 34.755 0.070 34.825 ;
    RECT 0 34.895 0.070 34.965 ;
    RECT 0 35.035 0.070 35.105 ;
    RECT 0 35.175 0.070 35.245 ;
    RECT 0 35.315 0.070 35.385 ;
    RECT 0 35.455 0.070 35.525 ;
    RECT 0 35.595 0.070 35.665 ;
    RECT 0 35.735 0.070 35.805 ;
    RECT 0 35.875 0.070 35.945 ;
    RECT 0 36.015 0.070 36.085 ;
    RECT 0 36.155 0.070 36.225 ;
    RECT 0 36.295 0.070 36.365 ;
    RECT 0 36.435 0.070 36.505 ;
    RECT 0 36.575 0.070 36.645 ;
    RECT 0 36.715 0.070 36.785 ;
    RECT 0 36.855 0.070 36.925 ;
    RECT 0 36.995 0.070 37.065 ;
    RECT 0 37.135 0.070 37.205 ;
    RECT 0 37.275 0.070 37.345 ;
    RECT 0 37.415 0.070 37.485 ;
    RECT 0 37.555 0.070 37.625 ;
    RECT 0 37.695 0.070 37.765 ;
    RECT 0 37.835 0.070 37.905 ;
    RECT 0 37.975 0.070 38.045 ;
    RECT 0 38.115 0.070 38.185 ;
    RECT 0 38.255 0.070 38.325 ;
    RECT 0 38.395 0.070 38.465 ;
    RECT 0 38.535 0.070 38.605 ;
    RECT 0 38.675 0.070 38.745 ;
    RECT 0 38.815 0.070 38.885 ;
    RECT 0 38.955 0.070 39.025 ;
    RECT 0 39.095 0.070 39.165 ;
    RECT 0 39.235 0.070 39.305 ;
    RECT 0 39.375 0.070 39.445 ;
    RECT 0 39.515 0.070 39.585 ;
    RECT 0 39.655 0.070 39.725 ;
    RECT 0 39.795 0.070 39.865 ;
    RECT 0 39.935 0.070 40.005 ;
    RECT 0 40.075 0.070 40.145 ;
    RECT 0 40.215 0.070 40.285 ;
    RECT 0 40.355 0.070 40.425 ;
    RECT 0 40.495 0.070 40.565 ;
    RECT 0 40.635 0.070 40.705 ;
    RECT 0 40.775 0.070 40.845 ;
    RECT 0 40.915 0.070 40.985 ;
    RECT 0 41.055 0.070 41.125 ;
    RECT 0 41.195 0.070 41.265 ;
    RECT 0 41.335 0.070 41.405 ;
    RECT 0 41.475 0.070 41.545 ;
    RECT 0 41.615 0.070 41.685 ;
    RECT 0 41.755 0.070 41.825 ;
    RECT 0 41.895 0.070 41.965 ;
    RECT 0 42.035 0.070 42.105 ;
    RECT 0 42.175 0.070 42.245 ;
    RECT 0 42.315 0.070 42.385 ;
    RECT 0 42.455 0.070 42.525 ;
    RECT 0 42.595 0.070 42.665 ;
    RECT 0 42.735 0.070 42.805 ;
    RECT 0 42.875 0.070 42.945 ;
    RECT 0 43.015 0.070 43.085 ;
    RECT 0 43.155 0.070 43.225 ;
    RECT 0 43.295 0.070 43.365 ;
    RECT 0 43.435 0.070 43.505 ;
    RECT 0 43.575 0.070 43.645 ;
    RECT 0 43.715 0.070 43.785 ;
    RECT 0 43.855 0.070 43.925 ;
    RECT 0 43.995 0.070 44.065 ;
    RECT 0 44.135 0.070 44.205 ;
    RECT 0 44.275 0.070 44.345 ;
    RECT 0 44.415 0.070 44.485 ;
    RECT 0 44.555 0.070 44.625 ;
    RECT 0 44.695 0.070 44.765 ;
    RECT 0 44.835 0.070 44.905 ;
    RECT 0 44.975 0.070 45.045 ;
    RECT 0 45.115 0.070 45.185 ;
    RECT 0 45.255 0.070 45.325 ;
    RECT 0 45.395 0.070 45.465 ;
    RECT 0 45.535 0.070 45.605 ;
    RECT 0 45.675 0.070 45.745 ;
    RECT 0 45.815 0.070 45.885 ;
    RECT 0 45.955 0.070 46.025 ;
    RECT 0 46.095 0.070 46.165 ;
    RECT 0 46.235 0.070 46.305 ;
    RECT 0 46.375 0.070 46.445 ;
    RECT 0 46.515 0.070 46.585 ;
    RECT 0 46.655 0.070 46.725 ;
    RECT 0 46.795 0.070 46.865 ;
    RECT 0 46.935 0.070 47.005 ;
    RECT 0 47.075 0.070 47.145 ;
    RECT 0 47.215 0.070 47.285 ;
    RECT 0 47.355 0.070 47.425 ;
    RECT 0 47.495 0.070 47.565 ;
    RECT 0 47.635 0.070 47.705 ;
    RECT 0 47.775 0.070 47.845 ;
    RECT 0 47.915 0.070 47.985 ;
    RECT 0 48.055 0.070 48.125 ;
    RECT 0 48.195 0.070 48.265 ;
    RECT 0 48.335 0.070 48.405 ;
    RECT 0 48.475 0.070 48.545 ;
    RECT 0 48.615 0.070 48.685 ;
    RECT 0 48.755 0.070 48.825 ;
    RECT 0 48.895 0.070 48.965 ;
    RECT 0 49.035 0.070 49.105 ;
    RECT 0 49.175 0.070 49.245 ;
    RECT 0 49.315 0.070 49.385 ;
    RECT 0 49.455 0.070 49.525 ;
    RECT 0 49.595 0.070 49.665 ;
    RECT 0 49.735 0.070 49.805 ;
    RECT 0 49.875 0.070 49.945 ;
    RECT 0 50.015 0.070 50.085 ;
    RECT 0 50.155 0.070 50.225 ;
    RECT 0 50.295 0.070 50.365 ;
    RECT 0 50.435 0.070 50.505 ;
    RECT 0 50.575 0.070 50.645 ;
    RECT 0 50.715 0.070 50.785 ;
    RECT 0 50.855 0.070 50.925 ;
    RECT 0 50.995 0.070 51.065 ;
    RECT 0 51.135 0.070 51.205 ;
    RECT 0 51.275 0.070 51.345 ;
    RECT 0 51.415 0.070 51.485 ;
    RECT 0 51.555 0.070 51.625 ;
    RECT 0 51.695 0.070 51.765 ;
    RECT 0 51.835 0.070 51.905 ;
    RECT 0 51.975 0.070 52.045 ;
    RECT 0 52.115 0.070 52.185 ;
    RECT 0 52.255 0.070 52.325 ;
    RECT 0 52.395 0.070 52.465 ;
    RECT 0 52.535 0.070 52.605 ;
    RECT 0 52.675 0.070 52.745 ;
    RECT 0 52.815 0.070 52.885 ;
    RECT 0 52.955 0.070 53.025 ;
    RECT 0 53.095 0.070 53.165 ;
    RECT 0 53.235 0.070 53.305 ;
    RECT 0 53.375 0.070 53.445 ;
    RECT 0 53.515 0.070 53.585 ;
    RECT 0 53.655 0.070 53.725 ;
    RECT 0 53.795 0.070 53.865 ;
    RECT 0 53.935 0.070 54.005 ;
    RECT 0 54.075 0.070 54.145 ;
    RECT 0 54.215 0.070 54.285 ;
    RECT 0 54.355 0.070 54.425 ;
    RECT 0 54.495 0.070 54.565 ;
    RECT 0 54.635 0.070 54.705 ;
    RECT 0 54.775 0.070 54.845 ;
    RECT 0 54.915 0.070 54.985 ;
    RECT 0 55.055 0.070 55.125 ;
    RECT 0 55.195 0.070 55.265 ;
    RECT 0 55.335 0.070 55.405 ;
    RECT 0 55.475 0.070 55.545 ;
    RECT 0 55.615 0.070 55.685 ;
    RECT 0 55.755 0.070 55.825 ;
    RECT 0 55.895 0.070 55.965 ;
    RECT 0 56.035 0.070 56.105 ;
    RECT 0 56.175 0.070 56.245 ;
    RECT 0 56.315 0.070 56.385 ;
    RECT 0 56.455 0.070 56.525 ;
    RECT 0 56.595 0.070 56.665 ;
    RECT 0 56.735 0.070 56.805 ;
    RECT 0 56.875 0.070 56.945 ;
    RECT 0 57.015 0.070 57.085 ;
    RECT 0 57.155 0.070 57.225 ;
    RECT 0 57.295 0.070 57.365 ;
    RECT 0 57.435 0.070 57.505 ;
    RECT 0 57.575 0.070 57.645 ;
    RECT 0 57.715 0.070 57.785 ;
    RECT 0 57.855 0.070 57.925 ;
    RECT 0 57.995 0.070 58.065 ;
    RECT 0 58.135 0.070 58.205 ;
    RECT 0 58.275 0.070 58.345 ;
    RECT 0 58.415 0.070 58.485 ;
    RECT 0 58.555 0.070 58.625 ;
    RECT 0 58.695 0.070 58.765 ;
    RECT 0 58.835 0.070 58.905 ;
    RECT 0 58.975 0.070 59.045 ;
    RECT 0 59.115 0.070 59.185 ;
    RECT 0 59.255 0.070 59.325 ;
    RECT 0 59.395 0.070 59.465 ;
    RECT 0 59.535 0.070 59.605 ;
    RECT 0 59.675 0.070 59.745 ;
    RECT 0 59.815 0.070 59.885 ;
    RECT 0 59.955 0.070 60.025 ;
    RECT 0 60.095 0.070 60.165 ;
    RECT 0 60.235 0.070 60.305 ;
    RECT 0 60.375 0.070 60.445 ;
    RECT 0 60.515 0.070 60.585 ;
    RECT 0 60.655 0.070 60.725 ;
    RECT 0 60.795 0.070 60.865 ;
    RECT 0 60.935 0.070 61.005 ;
    RECT 0 61.075 0.070 61.145 ;
    RECT 0 61.215 0.070 61.285 ;
    RECT 0 61.355 0.070 61.425 ;
    RECT 0 61.495 0.070 61.565 ;
    RECT 0 61.635 0.070 61.705 ;
    RECT 0 61.775 0.070 61.845 ;
    RECT 0 61.915 0.070 61.985 ;
    RECT 0 62.055 0.070 62.125 ;
    RECT 0 62.195 0.070 62.265 ;
    RECT 0 62.335 0.070 62.405 ;
    RECT 0 62.475 0.070 62.545 ;
    RECT 0 62.615 0.070 62.685 ;
    RECT 0 62.755 0.070 62.825 ;
    RECT 0 62.895 0.070 62.965 ;
    RECT 0 63.035 0.070 63.105 ;
    RECT 0 63.175 0.070 63.245 ;
    RECT 0 63.315 0.070 63.385 ;
    RECT 0 63.455 0.070 63.525 ;
    RECT 0 63.595 0.070 63.665 ;
    RECT 0 63.735 0.070 63.805 ;
    RECT 0 63.875 0.070 63.945 ;
    RECT 0 64.015 0.070 64.085 ;
    RECT 0 64.155 0.070 64.225 ;
    RECT 0 64.295 0.070 64.365 ;
    RECT 0 64.435 0.070 64.505 ;
    RECT 0 64.575 0.070 64.645 ;
    RECT 0 64.715 0.070 64.785 ;
    RECT 0 64.855 0.070 64.925 ;
    RECT 0 64.995 0.070 65.065 ;
    RECT 0 65.135 0.070 65.205 ;
    RECT 0 65.275 0.070 65.345 ;
    RECT 0 65.415 0.070 65.485 ;
    RECT 0 65.555 0.070 65.625 ;
    RECT 0 65.695 0.070 65.765 ;
    RECT 0 65.835 0.070 65.905 ;
    RECT 0 65.975 0.070 66.045 ;
    RECT 0 66.115 0.070 66.185 ;
    RECT 0 66.255 0.070 66.325 ;
    RECT 0 66.395 0.070 66.465 ;
    RECT 0 66.535 0.070 66.605 ;
    RECT 0 66.675 0.070 66.745 ;
    RECT 0 66.815 0.070 66.885 ;
    RECT 0 66.955 0.070 67.025 ;
    RECT 0 67.095 0.070 67.165 ;
    RECT 0 67.235 0.070 67.305 ;
    RECT 0 67.375 0.070 67.445 ;
    RECT 0 67.515 0.070 67.585 ;
    RECT 0 67.655 0.070 67.725 ;
    RECT 0 67.795 0.070 67.865 ;
    RECT 0 67.935 0.070 68.005 ;
    RECT 0 68.075 0.070 68.145 ;
    RECT 0 68.215 0.070 68.285 ;
    RECT 0 68.355 0.070 68.425 ;
    RECT 0 68.495 0.070 68.565 ;
    RECT 0 68.635 0.070 68.705 ;
    RECT 0 68.775 0.070 68.845 ;
    RECT 0 68.915 0.070 68.985 ;
    RECT 0 69.055 0.070 69.125 ;
    RECT 0 69.195 0.070 69.265 ;
    RECT 0 69.335 0.070 69.405 ;
    RECT 0 69.475 0.070 69.545 ;
    RECT 0 69.615 0.070 69.685 ;
    RECT 0 69.755 0.070 69.825 ;
    RECT 0 69.895 0.070 69.965 ;
    RECT 0 70.035 0.070 70.105 ;
    RECT 0 70.175 0.070 70.245 ;
    RECT 0 70.315 0.070 70.385 ;
    RECT 0 70.455 0.070 70.525 ;
    RECT 0 70.595 0.070 70.665 ;
    RECT 0 70.735 0.070 70.805 ;
    RECT 0 70.875 0.070 70.945 ;
    RECT 0 71.015 0.070 71.085 ;
    RECT 0 71.155 0.070 71.225 ;
    RECT 0 71.295 0.070 71.365 ;
    RECT 0 71.435 0.070 71.505 ;
    RECT 0 71.575 0.070 71.645 ;
    RECT 0 71.715 0.070 71.785 ;
    RECT 0 71.855 0.070 71.925 ;
    RECT 0 71.995 0.070 72.065 ;
    RECT 0 72.135 0.070 72.205 ;
    RECT 0 72.275 0.070 72.345 ;
    RECT 0 72.415 0.070 72.485 ;
    RECT 0 72.555 0.070 72.625 ;
    RECT 0 72.695 0.070 72.765 ;
    RECT 0 72.835 0.070 72.905 ;
    RECT 0 72.975 0.070 73.045 ;
    RECT 0 73.115 0.070 73.185 ;
    RECT 0 73.255 0.070 73.325 ;
    RECT 0 73.395 0.070 73.465 ;
    RECT 0 73.535 0.070 73.605 ;
    RECT 0 73.675 0.070 73.745 ;
    RECT 0 73.815 0.070 73.885 ;
    RECT 0 73.955 0.070 74.025 ;
    RECT 0 74.095 0.070 74.165 ;
    RECT 0 74.235 0.070 74.305 ;
    RECT 0 74.375 0.070 74.445 ;
    RECT 0 74.515 0.070 74.585 ;
    RECT 0 74.655 0.070 74.725 ;
    RECT 0 74.795 0.070 74.865 ;
    RECT 0 74.935 0.070 75.005 ;
    RECT 0 75.075 0.070 75.145 ;
    RECT 0 75.215 0.070 75.285 ;
    RECT 0 75.355 0.070 75.425 ;
    RECT 0 75.495 0.070 75.565 ;
    RECT 0 75.635 0.070 75.705 ;
    RECT 0 75.775 0.070 75.845 ;
    RECT 0 75.915 0.070 75.985 ;
    RECT 0 76.055 0.070 76.125 ;
    RECT 0 76.195 0.070 76.265 ;
    RECT 0 76.335 0.070 76.405 ;
    RECT 0 76.475 0.070 76.545 ;
    RECT 0 76.615 0.070 76.685 ;
    RECT 0 76.755 0.070 76.825 ;
    RECT 0 76.895 0.070 76.965 ;
    RECT 0 77.035 0.070 77.105 ;
    RECT 0 77.175 0.070 77.245 ;
    RECT 0 77.315 0.070 77.385 ;
    RECT 0 77.455 0.070 77.525 ;
    RECT 0 77.595 0.070 77.665 ;
    RECT 0 77.735 0.070 77.805 ;
    RECT 0 77.875 0.070 77.945 ;
    RECT 0 78.015 0.070 78.085 ;
    RECT 0 78.155 0.070 78.225 ;
    RECT 0 78.295 0.070 78.365 ;
    RECT 0 78.435 0.070 78.505 ;
    RECT 0 78.575 0.070 78.645 ;
    RECT 0 78.715 0.070 78.785 ;
    RECT 0 78.855 0.070 78.925 ;
    RECT 0 78.995 0.070 79.065 ;
    RECT 0 79.135 0.070 79.205 ;
    RECT 0 79.275 0.070 79.345 ;
    RECT 0 79.415 0.070 79.485 ;
    RECT 0 79.555 0.070 79.625 ;
    RECT 0 79.695 0.070 79.765 ;
    RECT 0 79.835 0.070 79.905 ;
    RECT 0 79.975 0.070 80.045 ;
    RECT 0 80.115 0.070 80.185 ;
    RECT 0 80.255 0.070 80.325 ;
    RECT 0 80.395 0.070 80.465 ;
    RECT 0 80.535 0.070 80.605 ;
    RECT 0 80.675 0.070 80.745 ;
    RECT 0 80.815 0.070 80.885 ;
    RECT 0 80.955 0.070 81.025 ;
    RECT 0 81.095 0.070 81.165 ;
    RECT 0 81.235 0.070 81.305 ;
    RECT 0 81.375 0.070 81.445 ;
    RECT 0 81.515 0.070 81.585 ;
    RECT 0 81.655 0.070 81.725 ;
    RECT 0 81.795 0.070 81.865 ;
    RECT 0 81.935 0.070 82.005 ;
    RECT 0 82.075 0.070 82.145 ;
    RECT 0 82.215 0.070 82.285 ;
    RECT 0 82.355 0.070 82.425 ;
    RECT 0 82.495 0.070 82.565 ;
    RECT 0 82.635 0.070 82.705 ;
    RECT 0 82.775 0.070 82.845 ;
    RECT 0 82.915 0.070 82.985 ;
    RECT 0 83.055 0.070 83.125 ;
    RECT 0 83.195 0.070 83.265 ;
    RECT 0 83.335 0.070 83.405 ;
    RECT 0 83.475 0.070 83.545 ;
    RECT 0 83.615 0.070 83.685 ;
    RECT 0 83.755 0.070 83.825 ;
    RECT 0 83.895 0.070 83.965 ;
    RECT 0 84.035 0.070 84.105 ;
    RECT 0 84.175 0.070 84.245 ;
    RECT 0 84.315 0.070 84.385 ;
    RECT 0 84.455 0.070 84.525 ;
    RECT 0 84.595 0.070 84.665 ;
    RECT 0 84.735 0.070 84.805 ;
    RECT 0 84.875 0.070 84.945 ;
    RECT 0 85.015 0.070 85.085 ;
    RECT 0 85.155 0.070 85.225 ;
    RECT 0 85.295 0.070 85.365 ;
    RECT 0 85.435 0.070 85.505 ;
    RECT 0 85.575 0.070 85.645 ;
    RECT 0 85.715 0.070 85.785 ;
    RECT 0 85.855 0.070 85.925 ;
    RECT 0 85.995 0.070 86.065 ;
    RECT 0 86.135 0.070 86.205 ;
    RECT 0 86.275 0.070 86.345 ;
    RECT 0 86.415 0.070 86.485 ;
    RECT 0 86.555 0.070 86.625 ;
    RECT 0 86.695 0.070 86.765 ;
    RECT 0 86.835 0.070 86.905 ;
    RECT 0 86.975 0.070 87.045 ;
    RECT 0 87.115 0.070 87.185 ;
    RECT 0 87.255 0.070 87.325 ;
    RECT 0 87.395 0.070 87.465 ;
    RECT 0 87.535 0.070 87.605 ;
    RECT 0 87.675 0.070 87.745 ;
    RECT 0 87.815 0.070 87.885 ;
    RECT 0 87.955 0.070 88.025 ;
    RECT 0 88.095 0.070 88.165 ;
    RECT 0 88.235 0.070 88.305 ;
    RECT 0 88.375 0.070 88.445 ;
    RECT 0 88.515 0.070 88.585 ;
    RECT 0 88.655 0.070 88.725 ;
    RECT 0 88.795 0.070 88.865 ;
    RECT 0 88.935 0.070 89.005 ;
    RECT 0 89.075 0.070 89.145 ;
    RECT 0 89.215 0.070 89.285 ;
    RECT 0 89.355 0.070 89.425 ;
    RECT 0 89.495 0.070 89.565 ;
    RECT 0 89.635 0.070 89.705 ;
    RECT 0 89.775 0.070 89.845 ;
    RECT 0 89.915 0.070 89.985 ;
    RECT 0 90.055 0.070 90.125 ;
    RECT 0 90.195 0.070 90.265 ;
    RECT 0 90.335 0.070 90.405 ;
    RECT 0 90.475 0.070 90.545 ;
    RECT 0 90.615 0.070 90.685 ;
    RECT 0 90.755 0.070 90.825 ;
    RECT 0 90.895 0.070 90.965 ;
    RECT 0 91.035 0.070 91.105 ;
    RECT 0 91.175 0.070 91.245 ;
    RECT 0 91.315 0.070 91.385 ;
    RECT 0 91.455 0.070 91.525 ;
    RECT 0 91.595 0.070 91.665 ;
    RECT 0 91.735 0.070 91.805 ;
    RECT 0 91.875 0.070 91.945 ;
    RECT 0 92.015 0.070 92.085 ;
    RECT 0 92.155 0.070 92.225 ;
    RECT 0 92.295 0.070 92.365 ;
    RECT 0 92.435 0.070 92.505 ;
    RECT 0 92.575 0.070 92.645 ;
    RECT 0 92.715 0.070 92.785 ;
    RECT 0 92.855 0.070 92.925 ;
    RECT 0 92.995 0.070 93.065 ;
    RECT 0 93.135 0.070 93.205 ;
    RECT 0 93.275 0.070 93.345 ;
    RECT 0 93.415 0.070 93.485 ;
    RECT 0 93.555 0.070 93.625 ;
    RECT 0 93.695 0.070 93.765 ;
    RECT 0 93.835 0.070 93.905 ;
    RECT 0 93.975 0.070 94.045 ;
    RECT 0 94.115 0.070 94.185 ;
    RECT 0 94.255 0.070 94.325 ;
    RECT 0 94.395 0.070 94.465 ;
    RECT 0 94.535 0.070 94.605 ;
    RECT 0 94.675 0.070 94.745 ;
    RECT 0 94.815 0.070 94.885 ;
    RECT 0 94.955 0.070 95.025 ;
    RECT 0 95.095 0.070 95.165 ;
    RECT 0 95.235 0.070 95.305 ;
    RECT 0 95.375 0.070 95.445 ;
    RECT 0 95.515 0.070 95.585 ;
    RECT 0 95.655 0.070 95.725 ;
    RECT 0 95.795 0.070 95.865 ;
    RECT 0 95.935 0.070 96.005 ;
    RECT 0 96.075 0.070 96.145 ;
    RECT 0 96.215 0.070 96.285 ;
    RECT 0 96.355 0.070 96.425 ;
    RECT 0 96.495 0.070 96.565 ;
    RECT 0 96.635 0.070 96.705 ;
    RECT 0 96.775 0.070 96.845 ;
    RECT 0 96.915 0.070 96.985 ;
    RECT 0 97.055 0.070 97.125 ;
    RECT 0 97.195 0.070 97.265 ;
    RECT 0 97.335 0.070 97.405 ;
    RECT 0 97.475 0.070 97.545 ;
    RECT 0 97.615 0.070 97.685 ;
    RECT 0 97.755 0.070 97.825 ;
    RECT 0 97.895 0.070 97.965 ;
    RECT 0 98.035 0.070 98.105 ;
    RECT 0 98.175 0.070 98.245 ;
    RECT 0 98.315 0.070 98.385 ;
    RECT 0 98.455 0.070 98.525 ;
    RECT 0 98.595 0.070 98.665 ;
    RECT 0 98.735 0.070 98.805 ;
    RECT 0 98.875 0.070 98.945 ;
    RECT 0 99.015 0.070 99.085 ;
    RECT 0 99.155 0.070 99.225 ;
    RECT 0 99.295 0.070 99.365 ;
    RECT 0 99.435 0.070 99.505 ;
    RECT 0 99.575 0.070 99.645 ;
    RECT 0 99.715 0.070 99.785 ;
    RECT 0 99.855 0.070 99.925 ;
    RECT 0 99.995 0.070 100.065 ;
    RECT 0 100.135 0.070 100.205 ;
    RECT 0 100.275 0.070 100.345 ;
    RECT 0 100.415 0.070 100.485 ;
    RECT 0 100.555 0.070 100.625 ;
    RECT 0 100.695 0.070 100.765 ;
    RECT 0 100.835 0.070 100.905 ;
    RECT 0 100.975 0.070 101.045 ;
    RECT 0 101.115 0.070 101.185 ;
    RECT 0 101.255 0.070 101.325 ;
    RECT 0 101.395 0.070 101.465 ;
    RECT 0 101.535 0.070 101.605 ;
    RECT 0 101.675 0.070 101.745 ;
    RECT 0 101.815 0.070 101.885 ;
    RECT 0 101.955 0.070 102.025 ;
    RECT 0 102.095 0.070 102.165 ;
    RECT 0 102.235 0.070 102.305 ;
    RECT 0 102.375 0.070 102.445 ;
    RECT 0 102.515 0.070 102.585 ;
    RECT 0 102.655 0.070 102.725 ;
    RECT 0 102.795 0.070 102.865 ;
    RECT 0 102.935 0.070 103.005 ;
    RECT 0 103.075 0.070 103.145 ;
    RECT 0 103.215 0.070 103.285 ;
    RECT 0 103.355 0.070 103.425 ;
    RECT 0 103.495 0.070 103.565 ;
    RECT 0 103.635 0.070 103.705 ;
    RECT 0 103.775 0.070 103.845 ;
    RECT 0 103.915 0.070 103.985 ;
    RECT 0 104.055 0.070 104.125 ;
    RECT 0 104.195 0.070 104.265 ;
    RECT 0 104.335 0.070 104.405 ;
    RECT 0 104.475 0.070 104.545 ;
    RECT 0 104.615 0.070 104.685 ;
    RECT 0 104.755 0.070 104.825 ;
    RECT 0 104.895 0.070 104.965 ;
    RECT 0 105.035 0.070 105.105 ;
    RECT 0 105.175 0.070 105.245 ;
    RECT 0 105.315 0.070 105.385 ;
    RECT 0 105.455 0.070 105.525 ;
    RECT 0 105.595 0.070 105.665 ;
    RECT 0 105.735 0.070 105.805 ;
    RECT 0 105.875 0.070 105.945 ;
    RECT 0 106.015 0.070 106.085 ;
    RECT 0 106.155 0.070 106.225 ;
    RECT 0 106.295 0.070 106.365 ;
    RECT 0 106.435 0.070 106.505 ;
    RECT 0 106.575 0.070 106.645 ;
    RECT 0 106.715 0.070 106.785 ;
    RECT 0 106.855 0.070 106.925 ;
    RECT 0 106.995 0.070 107.065 ;
    RECT 0 107.135 0.070 107.205 ;
    RECT 0 107.275 0.070 107.345 ;
    RECT 0 107.415 0.070 107.485 ;
    RECT 0 107.555 0.070 107.625 ;
    RECT 0 107.695 0.070 107.765 ;
    RECT 0 107.835 0.070 107.905 ;
    RECT 0 107.975 0.070 108.045 ;
    RECT 0 108.115 0.070 108.185 ;
    RECT 0 108.255 0.070 108.325 ;
    RECT 0 108.395 0.070 108.465 ;
    RECT 0 108.535 0.070 108.605 ;
    RECT 0 108.675 0.070 108.745 ;
    RECT 0 108.815 0.070 108.885 ;
    RECT 0 108.955 0.070 109.025 ;
    RECT 0 109.095 0.070 109.165 ;
    RECT 0 109.235 0.070 109.305 ;
    RECT 0 109.375 0.070 109.445 ;
    RECT 0 109.515 0.070 109.585 ;
    RECT 0 109.655 0.070 109.725 ;
    RECT 0 109.795 0.070 109.865 ;
    RECT 0 109.935 0.070 110.005 ;
    RECT 0 110.075 0.070 110.145 ;
    RECT 0 110.215 0.070 110.285 ;
    RECT 0 110.355 0.070 110.425 ;
    RECT 0 110.495 0.070 110.565 ;
    RECT 0 110.635 0.070 110.705 ;
    RECT 0 110.775 0.070 110.845 ;
    RECT 0 110.915 0.070 110.985 ;
    RECT 0 111.055 0.070 111.125 ;
    RECT 0 111.195 0.070 111.265 ;
    RECT 0 111.335 0.070 111.405 ;
    RECT 0 111.475 0.070 111.545 ;
    RECT 0 111.615 0.070 111.685 ;
    RECT 0 111.755 0.070 111.825 ;
    RECT 0 111.895 0.070 111.965 ;
    RECT 0 112.035 0.070 112.105 ;
    RECT 0 112.175 0.070 112.245 ;
    RECT 0 112.315 0.070 112.385 ;
    RECT 0 112.455 0.070 112.525 ;
    RECT 0 112.595 0.070 112.665 ;
    RECT 0 112.735 0.070 112.805 ;
    RECT 0 112.875 0.070 112.945 ;
    RECT 0 113.015 0.070 113.085 ;
    RECT 0 113.155 0.070 113.225 ;
    RECT 0 113.295 0.070 113.365 ;
    RECT 0 113.435 0.070 113.505 ;
    RECT 0 113.575 0.070 113.645 ;
    RECT 0 113.715 0.070 113.785 ;
    RECT 0 113.855 0.070 113.925 ;
    RECT 0 113.995 0.070 114.065 ;
    RECT 0 114.135 0.070 114.205 ;
    RECT 0 114.275 0.070 114.345 ;
    RECT 0 114.415 0.070 114.485 ;
    RECT 0 114.555 0.070 114.625 ;
    RECT 0 114.695 0.070 114.765 ;
    RECT 0 114.835 0.070 114.905 ;
    RECT 0 114.975 0.070 115.045 ;
    RECT 0 115.115 0.070 115.185 ;
    RECT 0 115.255 0.070 115.325 ;
    RECT 0 115.395 0.070 115.465 ;
    RECT 0 115.535 0.070 115.605 ;
    RECT 0 115.675 0.070 115.745 ;
    RECT 0 115.815 0.070 115.885 ;
    RECT 0 115.955 0.070 116.025 ;
    RECT 0 116.095 0.070 116.165 ;
    RECT 0 116.235 0.070 116.305 ;
    RECT 0 116.375 0.070 116.445 ;
    RECT 0 116.515 0.070 116.585 ;
    RECT 0 116.655 0.070 116.725 ;
    RECT 0 116.795 0.070 116.865 ;
    RECT 0 116.935 0.070 117.005 ;
    RECT 0 117.075 0.070 117.145 ;
    RECT 0 117.215 0.070 117.285 ;
    RECT 0 117.355 0.070 117.425 ;
    RECT 0 117.495 0.070 117.565 ;
    RECT 0 117.635 0.070 117.705 ;
    RECT 0 117.775 0.070 117.845 ;
    RECT 0 117.915 0.070 117.985 ;
    RECT 0 118.055 0.070 118.125 ;
    RECT 0 118.195 0.070 118.265 ;
    RECT 0 118.335 0.070 118.405 ;
    RECT 0 118.475 0.070 118.545 ;
    RECT 0 118.615 0.070 118.685 ;
    RECT 0 118.755 0.070 118.825 ;
    RECT 0 118.895 0.070 118.965 ;
    RECT 0 119.035 0.070 119.105 ;
    RECT 0 119.175 0.070 119.245 ;
    RECT 0 119.315 0.070 119.385 ;
    RECT 0 119.455 0.070 119.525 ;
    RECT 0 119.595 0.070 119.665 ;
    RECT 0 119.735 0.070 119.805 ;
    RECT 0 119.875 0.070 119.945 ;
    RECT 0 120.015 0.070 120.085 ;
    RECT 0 120.155 0.070 120.225 ;
    RECT 0 120.295 0.070 120.365 ;
    RECT 0 120.435 0.070 120.505 ;
    RECT 0 120.575 0.070 120.645 ;
    RECT 0 120.715 0.070 120.785 ;
    RECT 0 120.855 0.070 120.925 ;
    RECT 0 120.995 0.070 121.065 ;
    RECT 0 121.135 0.070 121.205 ;
    RECT 0 121.275 0.070 121.345 ;
    RECT 0 121.415 0.070 121.485 ;
    RECT 0 121.555 0.070 121.625 ;
    RECT 0 121.695 0.070 121.765 ;
    RECT 0 121.835 0.070 121.905 ;
    RECT 0 121.975 0.070 122.045 ;
    RECT 0 122.115 0.070 122.185 ;
    RECT 0 122.255 0.070 122.325 ;
    RECT 0 122.395 0.070 122.465 ;
    RECT 0 122.535 0.070 122.605 ;
    RECT 0 122.675 0.070 122.745 ;
    RECT 0 122.815 0.070 122.885 ;
    RECT 0 122.955 0.070 123.025 ;
    RECT 0 123.095 0.070 123.165 ;
    RECT 0 123.235 0.070 123.305 ;
    RECT 0 123.375 0.070 123.445 ;
    RECT 0 123.515 0.070 123.585 ;
    RECT 0 123.655 0.070 123.725 ;
    RECT 0 123.795 0.070 123.865 ;
    RECT 0 123.935 0.070 124.005 ;
    RECT 0 124.075 0.070 124.145 ;
    RECT 0 124.215 0.070 124.285 ;
    RECT 0 124.355 0.070 124.425 ;
    RECT 0 124.495 0.070 124.565 ;
    RECT 0 124.635 0.070 124.705 ;
    RECT 0 124.775 0.070 124.845 ;
    RECT 0 124.915 0.070 124.985 ;
    RECT 0 125.055 0.070 125.125 ;
    RECT 0 125.195 0.070 125.265 ;
    RECT 0 125.335 0.070 125.405 ;
    RECT 0 125.475 0.070 125.545 ;
    RECT 0 125.615 0.070 125.685 ;
    RECT 0 125.755 0.070 125.825 ;
    RECT 0 125.895 0.070 125.965 ;
    RECT 0 126.035 0.070 126.105 ;
    RECT 0 126.175 0.070 126.245 ;
    RECT 0 126.315 0.070 126.385 ;
    RECT 0 126.455 0.070 126.525 ;
    RECT 0 126.595 0.070 126.665 ;
    RECT 0 126.735 0.070 126.805 ;
    RECT 0 126.875 0.070 126.945 ;
    RECT 0 127.015 0.070 127.085 ;
    RECT 0 127.155 0.070 127.225 ;
    RECT 0 127.295 0.070 127.365 ;
    RECT 0 127.435 0.070 127.505 ;
    RECT 0 127.575 0.070 127.645 ;
    RECT 0 127.715 0.070 127.785 ;
    RECT 0 127.855 0.070 127.925 ;
    RECT 0 127.995 0.070 128.065 ;
    RECT 0 128.135 0.070 128.205 ;
    RECT 0 128.275 0.070 128.345 ;
    RECT 0 128.415 0.070 128.485 ;
    RECT 0 128.555 0.070 128.625 ;
    RECT 0 128.695 0.070 128.765 ;
    RECT 0 128.835 0.070 128.905 ;
    RECT 0 128.975 0.070 129.045 ;
    RECT 0 129.115 0.070 129.185 ;
    RECT 0 129.255 0.070 129.325 ;
    RECT 0 129.395 0.070 129.465 ;
    RECT 0 129.535 0.070 129.605 ;
    RECT 0 129.675 0.070 129.745 ;
    RECT 0 129.815 0.070 129.885 ;
    RECT 0 129.955 0.070 130.025 ;
    RECT 0 130.095 0.070 130.165 ;
    RECT 0 130.235 0.070 130.305 ;
    RECT 0 130.375 0.070 130.445 ;
    RECT 0 130.515 0.070 130.585 ;
    RECT 0 130.655 0.070 130.725 ;
    RECT 0 130.795 0.070 130.865 ;
    RECT 0 130.935 0.070 131.005 ;
    RECT 0 131.075 0.070 131.145 ;
    RECT 0 131.215 0.070 131.285 ;
    RECT 0 131.355 0.070 131.425 ;
    RECT 0 131.495 0.070 131.565 ;
    RECT 0 131.635 0.070 131.705 ;
    RECT 0 131.775 0.070 131.845 ;
    RECT 0 131.915 0.070 131.985 ;
    RECT 0 132.055 0.070 132.125 ;
    RECT 0 132.195 0.070 132.265 ;
    RECT 0 132.335 0.070 132.405 ;
    RECT 0 132.475 0.070 132.545 ;
    RECT 0 132.615 0.070 132.685 ;
    RECT 0 132.755 0.070 132.825 ;
    RECT 0 132.895 0.070 132.965 ;
    RECT 0 133.035 0.070 133.105 ;
    RECT 0 133.175 0.070 133.245 ;
    RECT 0 133.315 0.070 133.385 ;
    RECT 0 133.455 0.070 133.525 ;
    RECT 0 133.595 0.070 133.665 ;
    RECT 0 133.735 0.070 133.805 ;
    RECT 0 133.875 0.070 133.945 ;
    RECT 0 134.015 0.070 134.085 ;
    RECT 0 134.155 0.070 134.225 ;
    RECT 0 134.295 0.070 134.365 ;
    RECT 0 134.435 0.070 134.505 ;
    RECT 0 134.575 0.070 134.645 ;
    RECT 0 134.715 0.070 134.785 ;
    RECT 0 134.855 0.070 134.925 ;
    RECT 0 134.995 0.070 135.065 ;
    RECT 0 135.135 0.070 135.205 ;
    RECT 0 135.275 0.070 135.345 ;
    RECT 0 135.415 0.070 135.485 ;
    RECT 0 135.555 0.070 135.625 ;
    RECT 0 135.695 0.070 135.765 ;
    RECT 0 135.835 0.070 135.905 ;
    RECT 0 135.975 0.070 136.045 ;
    RECT 0 136.115 0.070 136.185 ;
    RECT 0 136.255 0.070 136.325 ;
    RECT 0 136.395 0.070 136.465 ;
    RECT 0 136.535 0.070 136.605 ;
    RECT 0 136.675 0.070 136.745 ;
    RECT 0 136.815 0.070 136.885 ;
    RECT 0 136.955 0.070 137.025 ;
    RECT 0 137.095 0.070 137.165 ;
    RECT 0 137.235 0.070 137.305 ;
    RECT 0 137.375 0.070 137.445 ;
    RECT 0 137.515 0.070 137.585 ;
    RECT 0 137.655 0.070 137.725 ;
    RECT 0 137.795 0.070 137.865 ;
    RECT 0 137.935 0.070 138.005 ;
    RECT 0 138.075 0.070 138.145 ;
    RECT 0 138.215 0.070 138.285 ;
    RECT 0 138.355 0.070 138.425 ;
    RECT 0 138.495 0.070 138.565 ;
    RECT 0 138.635 0.070 138.705 ;
    RECT 0 138.775 0.070 138.845 ;
    RECT 0 138.915 0.070 138.985 ;
    RECT 0 139.055 0.070 139.125 ;
    RECT 0 139.195 0.070 139.265 ;
    RECT 0 139.335 0.070 139.405 ;
    RECT 0 139.475 0.070 139.545 ;
    RECT 0 139.615 0.070 139.685 ;
    RECT 0 139.755 0.070 139.825 ;
    RECT 0 139.895 0.070 139.965 ;
    RECT 0 140.035 0.070 140.105 ;
    RECT 0 140.175 0.070 140.245 ;
    RECT 0 140.315 0.070 140.385 ;
    RECT 0 140.455 0.070 140.525 ;
    RECT 0 140.595 0.070 140.665 ;
    RECT 0 140.735 0.070 140.805 ;
    RECT 0 140.875 0.070 140.945 ;
    RECT 0 141.015 0.070 141.085 ;
    RECT 0 141.155 0.070 141.225 ;
    RECT 0 141.295 0.070 141.365 ;
    RECT 0 141.435 0.070 141.505 ;
    RECT 0 141.575 0.070 141.645 ;
    RECT 0 141.715 0.070 141.785 ;
    RECT 0 141.855 0.070 141.925 ;
    RECT 0 141.995 0.070 142.065 ;
    RECT 0 142.135 0.070 142.205 ;
    RECT 0 142.275 0.070 142.345 ;
    RECT 0 142.415 0.070 142.485 ;
    RECT 0 142.555 0.070 142.625 ;
    RECT 0 142.695 0.070 142.765 ;
    RECT 0 142.835 0.070 142.905 ;
    RECT 0 142.975 0.070 143.045 ;
    RECT 0 143.115 0.070 143.185 ;
    RECT 0 143.255 0.070 143.325 ;
    RECT 0 143.395 0.070 143.465 ;
    RECT 0 143.535 0.070 143.605 ;
    RECT 0 143.675 0.070 143.745 ;
    RECT 0 143.815 0.070 143.885 ;
    RECT 0 143.955 0.070 144.025 ;
    RECT 0 144.095 0.070 144.165 ;
    RECT 0 144.235 0.070 144.305 ;
    RECT 0 144.375 0.070 144.445 ;
    RECT 0 144.515 0.070 144.585 ;
    RECT 0 144.655 0.070 144.725 ;
    RECT 0 144.795 0.070 144.865 ;
    RECT 0 144.935 0.070 145.005 ;
    RECT 0 145.075 0.070 145.145 ;
    RECT 0 145.215 0.070 145.285 ;
    RECT 0 145.355 0.070 145.425 ;
    RECT 0 145.495 0.070 145.565 ;
    RECT 0 145.635 0.070 145.705 ;
    RECT 0 145.775 0.070 145.845 ;
    RECT 0 145.915 0.070 145.985 ;
    RECT 0 146.055 0.070 146.125 ;
    RECT 0 146.195 0.070 146.265 ;
    RECT 0 146.335 0.070 146.405 ;
    RECT 0 146.475 0.070 146.545 ;
    RECT 0 146.615 0.070 146.685 ;
    RECT 0 146.755 0.070 146.825 ;
    RECT 0 146.895 0.070 146.965 ;
    RECT 0 147.035 0.070 147.105 ;
    RECT 0 147.175 0.070 147.245 ;
    RECT 0 147.315 0.070 147.385 ;
    RECT 0 147.455 0.070 147.525 ;
    RECT 0 147.595 0.070 147.665 ;
    RECT 0 147.735 0.070 147.805 ;
    RECT 0 147.875 0.070 147.945 ;
    RECT 0 148.015 0.070 148.085 ;
    RECT 0 148.155 0.070 148.225 ;
    RECT 0 148.295 0.070 148.365 ;
    RECT 0 148.435 0.070 148.505 ;
    RECT 0 148.575 0.070 148.645 ;
    RECT 0 148.715 0.070 148.785 ;
    RECT 0 148.855 0.070 148.925 ;
    RECT 0 148.995 0.070 149.065 ;
    RECT 0 149.135 0.070 149.205 ;
    RECT 0 149.275 0.070 149.345 ;
    RECT 0 149.415 0.070 149.485 ;
    RECT 0 149.555 0.070 149.625 ;
    RECT 0 149.695 0.070 149.765 ;
    RECT 0 149.835 0.070 149.905 ;
    RECT 0 149.975 0.070 150.045 ;
    RECT 0 150.115 0.070 150.185 ;
    RECT 0 150.255 0.070 150.325 ;
    RECT 0 150.395 0.070 150.465 ;
    RECT 0 150.535 0.070 150.605 ;
    RECT 0 150.675 0.070 150.745 ;
    RECT 0 150.815 0.070 150.885 ;
    RECT 0 150.955 0.070 151.025 ;
    RECT 0 151.095 0.070 151.165 ;
    RECT 0 151.235 0.070 151.305 ;
    RECT 0 151.375 0.070 151.445 ;
    RECT 0 151.515 0.070 151.585 ;
    RECT 0 151.655 0.070 151.725 ;
    RECT 0 151.795 0.070 151.865 ;
    RECT 0 151.935 0.070 152.005 ;
    RECT 0 152.075 0.070 152.145 ;
    RECT 0 152.215 0.070 152.285 ;
    RECT 0 152.355 0.070 152.425 ;
    RECT 0 152.495 0.070 152.565 ;
    RECT 0 152.635 0.070 152.705 ;
    RECT 0 152.775 0.070 152.845 ;
    RECT 0 152.915 0.070 152.985 ;
    RECT 0 153.055 0.070 153.125 ;
    RECT 0 153.195 0.070 153.265 ;
    RECT 0 153.335 0.070 153.405 ;
    RECT 0 153.475 0.070 153.545 ;
    RECT 0 153.615 0.070 153.685 ;
    RECT 0 153.755 0.070 153.825 ;
    RECT 0 153.895 0.070 153.965 ;
    RECT 0 154.035 0.070 154.105 ;
    RECT 0 154.175 0.070 154.245 ;
    RECT 0 154.315 0.070 154.385 ;
    RECT 0 154.455 0.070 154.525 ;
    RECT 0 154.595 0.070 154.665 ;
    RECT 0 154.735 0.070 154.805 ;
    RECT 0 154.875 0.070 154.945 ;
    RECT 0 155.015 0.070 155.085 ;
    RECT 0 155.155 0.070 155.225 ;
    RECT 0 155.295 0.070 155.365 ;
    RECT 0 155.435 0.070 155.505 ;
    RECT 0 155.575 0.070 155.645 ;
    RECT 0 155.715 0.070 155.785 ;
    RECT 0 155.855 0.070 155.925 ;
    RECT 0 155.995 0.070 156.065 ;
    RECT 0 156.135 0.070 156.205 ;
    RECT 0 156.275 0.070 156.345 ;
    RECT 0 156.415 0.070 156.485 ;
    RECT 0 156.555 0.070 156.625 ;
    RECT 0 156.695 0.070 156.765 ;
    RECT 0 156.835 0.070 156.905 ;
    RECT 0 156.975 0.070 157.045 ;
    RECT 0 157.115 0.070 157.185 ;
    RECT 0 157.255 0.070 157.325 ;
    RECT 0 157.395 0.070 157.465 ;
    RECT 0 157.535 0.070 157.605 ;
    RECT 0 157.675 0.070 157.745 ;
    RECT 0 157.815 0.070 157.885 ;
    RECT 0 157.955 0.070 158.025 ;
    RECT 0 158.095 0.070 158.165 ;
    RECT 0 158.235 0.070 158.305 ;
    RECT 0 158.375 0.070 158.445 ;
    RECT 0 158.515 0.070 158.585 ;
    RECT 0 158.655 0.070 158.725 ;
    RECT 0 158.795 0.070 158.865 ;
    RECT 0 158.935 0.070 159.005 ;
    RECT 0 159.075 0.070 159.145 ;
    RECT 0 159.215 0.070 159.285 ;
    RECT 0 159.355 0.070 159.425 ;
    RECT 0 159.495 0.070 159.565 ;
    RECT 0 159.635 0.070 159.705 ;
    RECT 0 159.775 0.070 159.845 ;
    RECT 0 159.915 0.070 159.985 ;
    RECT 0 160.055 0.070 160.125 ;
    RECT 0 160.195 0.070 160.265 ;
    RECT 0 160.335 0.070 160.405 ;
    RECT 0 160.475 0.070 160.545 ;
    RECT 0 160.615 0.070 160.685 ;
    RECT 0 160.755 0.070 160.825 ;
    RECT 0 160.895 0.070 160.965 ;
    RECT 0 161.035 0.070 161.105 ;
    RECT 0 161.175 0.070 161.245 ;
    RECT 0 161.315 0.070 161.385 ;
    RECT 0 161.455 0.070 161.525 ;
    RECT 0 161.595 0.070 161.665 ;
    RECT 0 161.735 0.070 161.805 ;
    RECT 0 161.875 0.070 161.945 ;
    RECT 0 162.015 0.070 162.085 ;
    RECT 0 162.155 0.070 162.225 ;
    RECT 0 162.295 0.070 162.365 ;
    RECT 0 162.435 0.070 162.505 ;
    RECT 0 162.575 0.070 162.645 ;
    RECT 0 162.715 0.070 162.785 ;
    RECT 0 162.855 0.070 162.925 ;
    RECT 0 162.995 0.070 163.065 ;
    RECT 0 163.135 0.070 163.205 ;
    RECT 0 163.275 0.070 163.345 ;
    RECT 0 163.415 0.070 163.485 ;
    RECT 0 163.555 0.070 163.625 ;
    RECT 0 163.695 0.070 163.765 ;
    RECT 0 163.835 0.070 163.905 ;
    RECT 0 163.975 0.070 164.045 ;
    RECT 0 164.115 0.070 164.185 ;
    RECT 0 164.255 0.070 164.325 ;
    RECT 0 164.395 0.070 164.465 ;
    RECT 0 164.535 0.070 164.605 ;
    RECT 0 164.675 0.070 164.745 ;
    RECT 0 164.815 0.070 164.885 ;
    RECT 0 164.955 0.070 165.025 ;
    RECT 0 165.095 0.070 165.165 ;
    RECT 0 165.235 0.070 165.305 ;
    RECT 0 165.375 0.070 165.445 ;
    RECT 0 165.515 0.070 165.585 ;
    RECT 0 165.655 0.070 165.725 ;
    RECT 0 165.795 0.070 165.865 ;
    RECT 0 165.935 0.070 166.005 ;
    RECT 0 166.075 0.070 166.145 ;
    RECT 0 166.215 0.070 166.285 ;
    RECT 0 166.355 0.070 166.425 ;
    RECT 0 166.495 0.070 166.565 ;
    RECT 0 166.635 0.070 166.705 ;
    RECT 0 166.775 0.070 166.845 ;
    RECT 0 166.915 0.070 166.985 ;
    RECT 0 167.055 0.070 167.125 ;
    RECT 0 167.195 0.070 167.265 ;
    RECT 0 167.335 0.070 167.405 ;
    RECT 0 167.475 0.070 167.545 ;
    RECT 0 167.615 0.070 167.685 ;
    RECT 0 167.755 0.070 167.825 ;
    RECT 0 167.895 0.070 167.965 ;
    RECT 0 168.035 0.070 168.105 ;
    RECT 0 168.175 0.070 168.245 ;
    RECT 0 168.315 0.070 168.385 ;
    RECT 0 168.455 0.070 168.525 ;
    RECT 0 168.595 0.070 168.665 ;
    RECT 0 168.735 0.070 168.805 ;
    RECT 0 168.875 0.070 168.945 ;
    RECT 0 169.015 0.070 169.085 ;
    RECT 0 169.155 0.070 169.225 ;
    RECT 0 169.295 0.070 169.365 ;
    RECT 0 169.435 0.070 169.505 ;
    RECT 0 169.575 0.070 169.645 ;
    RECT 0 169.715 0.070 169.785 ;
    RECT 0 169.855 0.070 169.925 ;
    RECT 0 169.995 0.070 170.065 ;
    RECT 0 170.135 0.070 170.205 ;
    RECT 0 170.275 0.070 170.345 ;
    RECT 0 170.415 0.070 170.485 ;
    RECT 0 170.555 0.070 170.625 ;
    RECT 0 170.695 0.070 170.765 ;
    RECT 0 170.835 0.070 170.905 ;
    RECT 0 170.975 0.070 171.045 ;
    RECT 0 171.115 0.070 171.185 ;
    RECT 0 171.255 0.070 171.325 ;
    RECT 0 171.395 0.070 171.465 ;
    RECT 0 171.535 0.070 171.605 ;
    RECT 0 171.675 0.070 171.745 ;
    RECT 0 171.815 0.070 171.885 ;
    RECT 0 171.955 0.070 172.025 ;
    RECT 0 172.095 0.070 172.165 ;
    RECT 0 172.235 0.070 172.305 ;
    RECT 0 172.375 0.070 172.445 ;
    RECT 0 172.515 0.070 172.585 ;
    RECT 0 172.655 0.070 172.725 ;
    RECT 0 172.795 0.070 172.865 ;
    RECT 0 172.935 0.070 173.005 ;
    RECT 0 173.075 0.070 173.145 ;
    RECT 0 173.215 0.070 173.285 ;
    RECT 0 173.355 0.070 173.425 ;
    RECT 0 173.495 0.070 173.565 ;
    RECT 0 173.635 0.070 173.705 ;
    RECT 0 173.775 0.070 173.845 ;
    RECT 0 173.915 0.070 173.985 ;
    RECT 0 174.055 0.070 174.125 ;
    RECT 0 174.195 0.070 174.265 ;
    RECT 0 174.335 0.070 174.405 ;
    RECT 0 174.475 0.070 174.545 ;
    RECT 0 174.615 0.070 174.685 ;
    RECT 0 174.755 0.070 174.825 ;
    RECT 0 174.895 0.070 174.965 ;
    RECT 0 175.035 0.070 175.105 ;
    RECT 0 175.175 0.070 175.245 ;
    RECT 0 175.315 0.070 175.385 ;
    RECT 0 175.455 0.070 175.525 ;
    RECT 0 175.595 0.070 175.665 ;
    RECT 0 175.735 0.070 175.805 ;
    RECT 0 175.875 0.070 175.945 ;
    RECT 0 176.015 0.070 176.085 ;
    RECT 0 176.155 0.070 176.225 ;
    RECT 0 176.295 0.070 176.365 ;
    RECT 0 176.435 0.070 176.505 ;
    RECT 0 176.575 0.070 176.645 ;
    RECT 0 176.715 0.070 176.785 ;
    RECT 0 176.855 0.070 176.925 ;
    RECT 0 176.995 0.070 177.065 ;
    RECT 0 177.135 0.070 177.205 ;
    RECT 0 177.275 0.070 177.345 ;
    RECT 0 177.415 0.070 177.485 ;
    RECT 0 177.555 0.070 177.625 ;
    RECT 0 177.695 0.070 177.765 ;
    RECT 0 177.835 0.070 177.905 ;
    RECT 0 177.975 0.070 178.045 ;
    RECT 0 178.115 0.070 178.185 ;
    RECT 0 178.255 0.070 178.325 ;
    RECT 0 178.395 0.070 178.465 ;
    RECT 0 178.535 0.070 178.605 ;
    RECT 0 178.675 0.070 178.745 ;
    RECT 0 178.815 0.070 178.885 ;
    RECT 0 178.955 0.070 179.025 ;
    RECT 0 179.095 0.070 179.165 ;
    RECT 0 179.235 0.070 179.305 ;
    RECT 0 179.375 0.070 179.445 ;
    RECT 0 179.515 0.070 179.585 ;
    RECT 0 179.655 0.070 179.725 ;
    RECT 0 179.795 0.070 179.865 ;
    RECT 0 179.935 0.070 180.005 ;
    RECT 0 180.075 0.070 180.145 ;
    RECT 0 180.215 0.070 180.285 ;
    RECT 0 180.355 0.070 180.425 ;
    RECT 0 180.495 0.070 180.565 ;
    RECT 0 180.635 0.070 180.705 ;
    RECT 0 180.775 0.070 180.845 ;
    RECT 0 180.915 0.070 180.985 ;
    RECT 0 181.055 0.070 181.125 ;
    RECT 0 181.195 0.070 181.265 ;
    RECT 0 181.335 0.070 181.405 ;
    RECT 0 181.475 0.070 181.545 ;
    RECT 0 181.615 0.070 181.685 ;
    RECT 0 181.755 0.070 181.825 ;
    RECT 0 181.895 0.070 181.965 ;
    RECT 0 182.035 0.070 182.105 ;
    RECT 0 182.175 0.070 182.245 ;
    RECT 0 182.315 0.070 182.385 ;
    RECT 0 182.455 0.070 182.525 ;
    RECT 0 182.595 0.070 182.665 ;
    RECT 0 182.735 0.070 182.805 ;
    RECT 0 182.875 0.070 182.945 ;
    RECT 0 183.015 0.070 183.085 ;
    RECT 0 183.155 0.070 183.225 ;
    RECT 0 183.295 0.070 183.365 ;
    RECT 0 183.435 0.070 183.505 ;
    RECT 0 183.575 0.070 183.645 ;
    RECT 0 183.715 0.070 183.785 ;
    RECT 0 183.855 0.070 183.925 ;
    RECT 0 183.995 0.070 184.065 ;
    RECT 0 184.135 0.070 184.205 ;
    RECT 0 184.275 0.070 184.345 ;
    RECT 0 184.415 0.070 184.485 ;
    RECT 0 184.555 0.070 184.625 ;
    RECT 0 184.695 0.070 184.765 ;
    RECT 0 184.835 0.070 184.905 ;
    RECT 0 184.975 0.070 185.045 ;
    RECT 0 185.115 0.070 185.185 ;
    RECT 0 185.255 0.070 185.325 ;
    RECT 0 185.395 0.070 185.465 ;
    RECT 0 185.535 0.070 185.605 ;
    RECT 0 185.675 0.070 185.745 ;
    RECT 0 185.815 0.070 185.885 ;
    RECT 0 185.955 0.070 186.025 ;
    RECT 0 186.095 0.070 186.165 ;
    RECT 0 186.235 0.070 186.305 ;
    RECT 0 186.375 0.070 186.445 ;
    RECT 0 186.515 0.070 186.585 ;
    RECT 0 186.655 0.070 186.725 ;
    RECT 0 186.795 0.070 186.865 ;
    RECT 0 186.935 0.070 187.005 ;
    RECT 0 187.075 0.070 187.145 ;
    RECT 0 187.215 0.070 187.285 ;
    RECT 0 187.355 0.070 187.425 ;
    RECT 0 187.495 0.070 187.565 ;
    RECT 0 187.635 0.070 187.705 ;
    RECT 0 187.775 0.070 187.845 ;
    RECT 0 187.915 0.070 187.985 ;
    RECT 0 188.055 0.070 188.125 ;
    RECT 0 188.195 0.070 188.265 ;
    RECT 0 188.335 0.070 188.405 ;
    RECT 0 188.475 0.070 188.545 ;
    RECT 0 188.615 0.070 188.685 ;
    RECT 0 188.755 0.070 188.825 ;
    RECT 0 188.895 0.070 188.965 ;
    RECT 0 189.035 0.070 189.105 ;
    RECT 0 189.175 0.070 189.245 ;
    RECT 0 189.315 0.070 189.385 ;
    RECT 0 189.455 0.070 189.525 ;
    RECT 0 189.595 0.070 189.665 ;
    RECT 0 189.735 0.070 189.805 ;
    RECT 0 189.875 0.070 189.945 ;
    RECT 0 190.015 0.070 190.085 ;
    RECT 0 190.155 0.070 190.225 ;
    RECT 0 190.295 0.070 190.365 ;
    RECT 0 190.435 0.070 190.505 ;
    RECT 0 190.575 0.070 190.645 ;
    RECT 0 190.715 0.070 190.785 ;
    RECT 0 190.855 0.070 190.925 ;
    RECT 0 190.995 0.070 191.065 ;
    RECT 0 191.135 0.070 191.205 ;
    RECT 0 191.275 0.070 191.345 ;
    RECT 0 191.415 0.070 191.485 ;
    RECT 0 191.555 0.070 191.625 ;
    RECT 0 191.695 0.070 191.765 ;
    RECT 0 191.835 0.070 191.905 ;
    RECT 0 191.975 0.070 192.045 ;
    RECT 0 192.115 0.070 192.185 ;
    RECT 0 192.255 0.070 192.325 ;
    RECT 0 192.395 0.070 192.465 ;
    RECT 0 192.535 0.070 192.605 ;
    RECT 0 192.675 0.070 192.745 ;
    RECT 0 192.815 0.070 192.885 ;
    RECT 0 192.955 0.070 193.025 ;
    RECT 0 193.095 0.070 193.165 ;
    RECT 0 193.235 0.070 193.305 ;
    RECT 0 193.375 0.070 193.445 ;
    RECT 0 193.515 0.070 193.585 ;
    RECT 0 193.655 0.070 193.725 ;
    RECT 0 193.795 0.070 193.865 ;
    RECT 0 193.935 0.070 194.005 ;
    RECT 0 194.075 0.070 194.145 ;
    RECT 0 194.215 0.070 194.285 ;
    RECT 0 194.355 0.070 194.425 ;
    RECT 0 194.495 0.070 194.565 ;
    RECT 0 194.635 0.070 194.705 ;
    RECT 0 194.775 0.070 194.845 ;
    RECT 0 194.915 0.070 194.985 ;
    RECT 0 195.055 0.070 195.125 ;
    RECT 0 195.195 0.070 195.265 ;
    RECT 0 195.335 0.070 195.405 ;
    RECT 0 195.475 0.070 195.545 ;
    RECT 0 195.615 0.070 195.685 ;
    RECT 0 195.755 0.070 195.825 ;
    RECT 0 195.895 0.070 195.965 ;
    RECT 0 196.035 0.070 196.105 ;
    RECT 0 196.175 0.070 196.245 ;
    RECT 0 196.315 0.070 196.385 ;
    RECT 0 196.455 0.070 196.525 ;
    RECT 0 196.595 0.070 196.665 ;
    RECT 0 196.735 0.070 196.805 ;
    RECT 0 196.875 0.070 196.945 ;
    RECT 0 197.015 0.070 197.085 ;
    RECT 0 197.155 0.070 197.225 ;
    RECT 0 197.295 0.070 197.365 ;
    RECT 0 197.435 0.070 197.505 ;
    RECT 0 197.575 0.070 197.645 ;
    RECT 0 197.715 0.070 197.785 ;
    RECT 0 197.855 0.070 197.925 ;
    RECT 0 197.995 0.070 198.065 ;
    RECT 0 198.135 0.070 198.205 ;
    RECT 0 198.275 0.070 198.345 ;
    RECT 0 198.415 0.070 198.485 ;
    RECT 0 198.555 0.070 198.625 ;
    RECT 0 198.695 0.070 198.765 ;
    RECT 0 198.835 0.070 198.905 ;
    RECT 0 198.975 0.070 199.045 ;
    RECT 0 199.115 0.070 199.185 ;
    RECT 0 199.255 0.070 199.325 ;
    RECT 0 199.395 0.070 199.465 ;
    RECT 0 199.535 0.070 199.605 ;
    RECT 0 199.675 0.070 199.745 ;
    RECT 0 199.815 0.070 199.885 ;
    RECT 0 199.955 0.070 200.025 ;
    RECT 0 200.095 0.070 200.165 ;
    RECT 0 200.235 0.070 200.305 ;
    RECT 0 200.375 0.070 200.445 ;
    RECT 0 200.515 0.070 200.585 ;
    RECT 0 200.655 0.070 200.725 ;
    RECT 0 200.795 0.070 200.865 ;
    RECT 0 200.935 0.070 201.005 ;
    RECT 0 201.075 0.070 201.145 ;
    RECT 0 201.215 0.070 201.285 ;
    RECT 0 201.355 0.070 201.425 ;
    RECT 0 201.495 0.070 201.565 ;
    RECT 0 201.635 0.070 201.705 ;
    RECT 0 201.775 0.070 201.845 ;
    RECT 0 201.915 0.070 201.985 ;
    RECT 0 202.055 0.070 202.125 ;
    RECT 0 202.195 0.070 202.265 ;
    RECT 0 202.335 0.070 202.405 ;
    RECT 0 202.475 0.070 202.545 ;
    RECT 0 202.615 0.070 202.685 ;
    RECT 0 202.755 0.070 202.825 ;
    RECT 0 202.895 0.070 202.965 ;
    RECT 0 203.035 0.070 203.105 ;
    RECT 0 203.175 0.070 203.245 ;
    RECT 0 203.315 0.070 203.385 ;
    RECT 0 203.455 0.070 203.525 ;
    RECT 0 203.595 0.070 203.665 ;
    RECT 0 203.735 0.070 203.805 ;
    RECT 0 203.875 0.070 203.945 ;
    RECT 0 204.015 0.070 204.085 ;
    RECT 0 204.155 0.070 204.225 ;
    RECT 0 204.295 0.070 204.365 ;
    RECT 0 204.435 0.070 204.505 ;
    RECT 0 204.575 0.070 204.645 ;
    RECT 0 204.715 0.070 204.785 ;
    RECT 0 204.855 0.070 204.925 ;
    RECT 0 204.995 0.070 205.065 ;
    RECT 0 205.135 0.070 205.205 ;
    RECT 0 205.275 0.070 205.345 ;
    RECT 0 205.415 0.070 205.485 ;
    RECT 0 205.555 0.070 205.625 ;
    RECT 0 205.695 0.070 205.765 ;
    RECT 0 205.835 0.070 205.905 ;
    RECT 0 205.975 0.070 206.045 ;
    RECT 0 206.115 0.070 206.185 ;
    RECT 0 206.255 0.070 206.325 ;
    RECT 0 206.395 0.070 206.465 ;
    RECT 0 206.535 0.070 206.605 ;
    RECT 0 206.675 0.070 206.745 ;
    RECT 0 206.815 0.070 206.885 ;
    RECT 0 206.955 0.070 207.025 ;
    RECT 0 207.095 0.070 207.165 ;
    RECT 0 207.235 0.070 207.305 ;
    RECT 0 207.375 0.070 207.445 ;
    RECT 0 207.515 0.070 207.585 ;
    RECT 0 207.655 0.070 207.725 ;
    RECT 0 207.795 0.070 207.865 ;
    RECT 0 207.935 0.070 208.005 ;
    RECT 0 208.075 0.070 208.145 ;
    RECT 0 208.215 0.070 208.285 ;
    RECT 0 208.355 0.070 208.425 ;
    RECT 0 208.495 0.070 208.565 ;
    RECT 0 208.635 0.070 208.705 ;
    RECT 0 208.775 0.070 208.845 ;
    RECT 0 208.915 0.070 208.985 ;
    RECT 0 209.055 0.070 209.125 ;
    RECT 0 209.195 0.070 209.265 ;
    RECT 0 209.335 0.070 209.405 ;
    RECT 0 209.475 0.070 209.545 ;
    RECT 0 209.615 0.070 209.685 ;
    RECT 0 209.755 0.070 209.825 ;
    RECT 0 209.895 0.070 209.965 ;
    RECT 0 210.035 0.070 210.105 ;
    RECT 0 210.175 0.070 210.245 ;
    RECT 0 210.315 0.070 210.385 ;
    RECT 0 210.455 0.070 210.525 ;
    RECT 0 210.595 0.070 210.665 ;
    RECT 0 210.735 0.070 210.805 ;
    RECT 0 210.875 0.070 210.945 ;
    RECT 0 211.015 0.070 211.085 ;
    RECT 0 211.155 0.070 211.225 ;
    RECT 0 211.295 0.070 211.365 ;
    RECT 0 211.435 0.070 211.505 ;
    RECT 0 211.575 0.070 211.645 ;
    RECT 0 211.715 0.070 211.785 ;
    RECT 0 211.855 0.070 211.925 ;
    RECT 0 211.995 0.070 212.065 ;
    RECT 0 212.135 0.070 212.205 ;
    RECT 0 212.275 0.070 212.345 ;
    RECT 0 212.415 0.070 212.485 ;
    RECT 0 212.555 0.070 212.625 ;
    RECT 0 212.695 0.070 212.765 ;
    RECT 0 212.835 0.070 212.905 ;
    RECT 0 212.975 0.070 213.045 ;
    RECT 0 213.115 0.070 213.185 ;
    RECT 0 213.255 0.070 213.325 ;
    RECT 0 213.395 0.070 213.465 ;
    RECT 0 213.535 0.070 213.605 ;
    RECT 0 213.675 0.070 213.745 ;
    RECT 0 213.815 0.070 213.885 ;
    RECT 0 213.955 0.070 214.025 ;
    RECT 0 214.095 0.070 214.165 ;
    RECT 0 214.235 0.070 214.305 ;
    RECT 0 214.375 0.070 214.445 ;
    RECT 0 214.515 0.070 214.585 ;
    RECT 0 214.655 0.070 214.725 ;
    RECT 0 214.795 0.070 214.865 ;
    RECT 0 214.935 0.070 215.005 ;
    RECT 0 215.075 0.070 215.145 ;
    RECT 0 215.215 0.070 215.285 ;
    RECT 0 215.355 0.070 215.425 ;
    RECT 0 215.495 0.070 215.565 ;
    RECT 0 215.635 0.070 215.705 ;
    RECT 0 215.775 0.070 215.845 ;
    RECT 0 215.915 0.070 215.985 ;
    RECT 0 216.055 0.070 216.125 ;
    RECT 0 216.195 0.070 216.265 ;
    RECT 0 216.335 0.070 216.405 ;
    RECT 0 216.475 0.070 216.545 ;
    RECT 0 216.615 0.070 216.685 ;
    RECT 0 216.755 0.070 216.825 ;
    RECT 0 216.895 0.070 216.965 ;
    RECT 0 217.035 0.070 217.105 ;
    RECT 0 217.175 0.070 217.245 ;
    RECT 0 217.315 0.070 217.385 ;
    RECT 0 217.455 0.070 217.525 ;
    RECT 0 217.595 0.070 217.665 ;
    RECT 0 217.735 0.070 217.805 ;
    RECT 0 217.875 0.070 217.945 ;
    RECT 0 218.015 0.070 218.085 ;
    RECT 0 218.155 0.070 218.225 ;
    RECT 0 218.295 0.070 218.365 ;
    RECT 0 218.435 0.070 218.505 ;
    RECT 0 218.575 0.070 218.645 ;
    RECT 0 218.715 0.070 218.785 ;
    RECT 0 218.855 0.070 218.925 ;
    RECT 0 218.995 0.070 219.065 ;
    RECT 0 219.135 0.070 219.205 ;
    RECT 0 219.275 0.070 219.345 ;
    RECT 0 219.415 0.070 219.485 ;
    RECT 0 219.555 0.070 219.625 ;
    RECT 0 219.695 0.070 219.765 ;
    RECT 0 219.835 0.070 219.905 ;
    RECT 0 219.975 0.070 220.045 ;
    RECT 0 220.115 0.070 220.185 ;
    RECT 0 220.255 0.070 220.325 ;
    RECT 0 220.395 0.070 220.465 ;
    RECT 0 220.535 0.070 220.605 ;
    RECT 0 220.675 0.070 220.745 ;
    RECT 0 220.815 0.070 220.885 ;
    RECT 0 220.955 0.070 221.025 ;
    RECT 0 221.095 0.070 221.165 ;
    RECT 0 221.235 0.070 221.305 ;
    RECT 0 221.375 0.070 221.445 ;
    RECT 0 221.515 0.070 221.585 ;
    RECT 0 221.655 0.070 221.725 ;
    RECT 0 221.795 0.070 221.865 ;
    RECT 0 221.935 0.070 222.005 ;
    RECT 0 222.075 0.070 222.145 ;
    RECT 0 222.215 0.070 222.285 ;
    RECT 0 222.355 0.070 222.425 ;
    RECT 0 222.495 0.070 222.565 ;
    RECT 0 222.635 0.070 222.705 ;
    RECT 0 222.775 0.070 222.845 ;
    RECT 0 222.915 0.070 222.985 ;
    RECT 0 223.055 0.070 223.125 ;
    RECT 0 223.195 0.070 223.265 ;
    RECT 0 223.335 0.070 223.405 ;
    RECT 0 223.475 0.070 223.545 ;
    RECT 0 223.615 0.070 223.685 ;
    RECT 0 223.755 0.070 223.825 ;
    RECT 0 223.895 0.070 223.965 ;
    RECT 0 224.035 0.070 224.105 ;
    RECT 0 224.175 0.070 224.245 ;
    RECT 0 224.315 0.070 224.385 ;
    RECT 0 224.455 0.070 224.525 ;
    RECT 0 224.595 0.070 224.665 ;
    RECT 0 224.735 0.070 224.805 ;
    RECT 0 224.875 0.070 224.945 ;
    RECT 0 225.015 0.070 225.085 ;
    RECT 0 225.155 0.070 225.225 ;
    RECT 0 225.295 0.070 225.365 ;
    RECT 0 225.435 0.070 225.505 ;
    RECT 0 225.575 0.070 225.645 ;
    RECT 0 225.715 0.070 225.785 ;
    RECT 0 225.855 0.070 225.925 ;
    RECT 0 225.995 0.070 226.065 ;
    RECT 0 226.135 0.070 226.205 ;
    RECT 0 226.275 0.070 226.345 ;
    RECT 0 226.415 0.070 226.485 ;
    RECT 0 226.555 0.070 226.625 ;
    RECT 0 226.695 0.070 226.765 ;
    RECT 0 226.835 0.070 226.905 ;
    RECT 0 226.975 0.070 227.045 ;
    RECT 0 227.115 0.070 227.185 ;
    RECT 0 227.255 0.070 227.325 ;
    RECT 0 227.395 0.070 227.465 ;
    RECT 0 227.535 0.070 227.605 ;
    RECT 0 227.675 0.070 227.745 ;
    RECT 0 227.815 0.070 227.885 ;
    RECT 0 227.955 0.070 228.025 ;
    RECT 0 228.095 0.070 228.165 ;
    RECT 0 228.235 0.070 228.305 ;
    RECT 0 228.375 0.070 228.445 ;
    RECT 0 228.515 0.070 228.585 ;
    RECT 0 228.655 0.070 228.725 ;
    RECT 0 228.795 0.070 228.865 ;
    RECT 0 228.935 0.070 229.005 ;
    RECT 0 229.075 0.070 229.145 ;
    RECT 0 229.215 0.070 229.285 ;
    RECT 0 229.355 0.070 229.425 ;
    RECT 0 229.495 0.070 229.565 ;
    RECT 0 229.635 0.070 229.705 ;
    RECT 0 229.775 0.070 229.845 ;
    RECT 0 229.915 0.070 229.985 ;
    RECT 0 230.055 0.070 230.125 ;
    RECT 0 230.195 0.070 230.265 ;
    RECT 0 230.335 0.070 230.405 ;
    RECT 0 230.475 0.070 230.545 ;
    RECT 0 230.615 0.070 230.685 ;
    RECT 0 230.755 0.070 230.825 ;
    RECT 0 230.895 0.070 230.965 ;
    RECT 0 231.035 0.070 231.105 ;
    RECT 0 231.175 0.070 231.245 ;
    RECT 0 231.315 0.070 231.385 ;
    RECT 0 231.455 0.070 231.525 ;
    RECT 0 231.595 0.070 231.665 ;
    RECT 0 231.735 0.070 231.805 ;
    RECT 0 231.875 0.070 231.945 ;
    RECT 0 232.015 0.070 232.085 ;
    RECT 0 232.155 0.070 232.225 ;
    RECT 0 232.295 0.070 232.365 ;
    RECT 0 232.435 0.070 232.505 ;
    RECT 0 232.575 0.070 232.645 ;
    RECT 0 232.715 0.070 232.785 ;
    RECT 0 232.855 0.070 232.925 ;
    RECT 0 232.995 0.070 233.065 ;
    RECT 0 233.135 0.070 233.205 ;
    RECT 0 233.275 0.070 233.345 ;
    RECT 0 233.415 0.070 233.485 ;
    RECT 0 233.555 0.070 233.625 ;
    RECT 0 233.695 0.070 233.765 ;
    RECT 0 233.835 0.070 233.905 ;
    RECT 0 233.975 0.070 234.045 ;
    RECT 0 234.115 0.070 234.185 ;
    RECT 0 234.255 0.070 234.325 ;
    RECT 0 234.395 0.070 234.465 ;
    RECT 0 234.535 0.070 234.605 ;
    RECT 0 234.675 0.070 234.745 ;
    RECT 0 234.815 0.070 234.885 ;
    RECT 0 234.955 0.070 235.025 ;
    RECT 0 235.095 0.070 235.165 ;
    RECT 0 235.235 0.070 235.305 ;
    RECT 0 235.375 0.070 235.445 ;
    RECT 0 235.515 0.070 235.585 ;
    RECT 0 235.655 0.070 235.725 ;
    RECT 0 235.795 0.070 235.865 ;
    RECT 0 235.935 0.070 236.005 ;
    RECT 0 236.075 0.070 236.145 ;
    RECT 0 236.215 0.070 236.285 ;
    RECT 0 236.355 0.070 236.425 ;
    RECT 0 236.495 0.070 236.565 ;
    RECT 0 236.635 0.070 236.705 ;
    RECT 0 236.775 0.070 236.845 ;
    RECT 0 236.915 0.070 236.985 ;
    RECT 0 237.055 0.070 237.125 ;
    RECT 0 237.195 0.070 237.265 ;
    RECT 0 237.335 0.070 237.405 ;
    RECT 0 237.475 0.070 237.545 ;
    RECT 0 237.615 0.070 237.685 ;
    RECT 0 237.755 0.070 237.825 ;
    RECT 0 237.895 0.070 237.965 ;
    RECT 0 238.035 0.070 238.105 ;
    RECT 0 238.175 0.070 238.245 ;
    RECT 0 238.315 0.070 238.385 ;
    RECT 0 238.455 0.070 238.525 ;
    RECT 0 238.595 0.070 238.665 ;
    RECT 0 238.735 0.070 238.805 ;
    RECT 0 238.875 0.070 238.945 ;
    RECT 0 239.015 0.070 239.085 ;
    RECT 0 239.155 0.070 239.225 ;
    RECT 0 239.295 0.070 239.365 ;
    RECT 0 239.435 0.070 239.505 ;
    RECT 0 239.575 0.070 239.645 ;
    RECT 0 239.715 0.070 239.785 ;
    RECT 0 239.855 0.070 239.925 ;
    RECT 0 239.995 0.070 240.065 ;
    RECT 0 240.135 0.070 240.205 ;
    RECT 0 240.275 0.070 240.345 ;
    RECT 0 240.415 0.070 240.485 ;
    RECT 0 240.555 0.070 240.625 ;
    RECT 0 240.695 0.070 240.765 ;
    RECT 0 240.835 0.070 240.905 ;
    RECT 0 240.975 0.070 241.045 ;
    RECT 0 241.115 0.070 241.185 ;
    RECT 0 241.255 0.070 241.325 ;
    RECT 0 241.395 0.070 241.465 ;
    RECT 0 241.535 0.070 241.605 ;
    RECT 0 241.675 0.070 241.745 ;
    RECT 0 241.815 0.070 241.885 ;
    RECT 0 241.955 0.070 242.025 ;
    RECT 0 242.095 0.070 242.165 ;
    RECT 0 242.235 0.070 242.305 ;
    RECT 0 242.375 0.070 242.445 ;
    RECT 0 242.515 0.070 242.585 ;
    RECT 0 242.655 0.070 242.725 ;
    RECT 0 242.795 0.070 242.865 ;
    RECT 0 242.935 0.070 243.005 ;
    RECT 0 243.075 0.070 243.145 ;
    RECT 0 243.215 0.070 243.285 ;
    RECT 0 243.355 0.070 243.425 ;
    RECT 0 243.495 0.070 243.565 ;
    RECT 0 243.635 0.070 243.705 ;
    RECT 0 243.775 0.070 243.845 ;
    RECT 0 243.915 0.070 243.985 ;
    RECT 0 244.055 0.070 244.125 ;
    RECT 0 244.195 0.070 244.265 ;
    RECT 0 244.335 0.070 244.405 ;
    RECT 0 244.475 0.070 244.545 ;
    RECT 0 244.615 0.070 244.685 ;
    RECT 0 244.755 0.070 244.825 ;
    RECT 0 244.895 0.070 244.965 ;
    RECT 0 245.035 0.070 245.105 ;
    RECT 0 245.175 0.070 245.245 ;
    RECT 0 245.315 0.070 245.385 ;
    RECT 0 245.455 0.070 245.525 ;
    RECT 0 245.595 0.070 245.665 ;
    RECT 0 245.735 0.070 245.805 ;
    RECT 0 245.875 0.070 245.945 ;
    RECT 0 246.015 0.070 246.085 ;
    RECT 0 246.155 0.070 246.225 ;
    RECT 0 246.295 0.070 246.365 ;
    RECT 0 246.435 0.070 246.505 ;
    RECT 0 246.575 0.070 246.645 ;
    RECT 0 246.715 0.070 246.785 ;
    RECT 0 246.855 0.070 246.925 ;
    RECT 0 246.995 0.070 247.065 ;
    RECT 0 247.135 0.070 247.205 ;
    RECT 0 247.275 0.070 247.345 ;
    RECT 0 247.415 0.070 247.485 ;
    RECT 0 247.555 0.070 247.625 ;
    RECT 0 247.695 0.070 247.765 ;
    RECT 0 247.835 0.070 247.905 ;
    RECT 0 247.975 0.070 248.045 ;
    RECT 0 248.115 0.070 248.185 ;
    RECT 0 248.255 0.070 248.325 ;
    RECT 0 248.395 0.070 248.465 ;
    RECT 0 248.535 0.070 248.605 ;
    RECT 0 248.675 0.070 248.745 ;
    RECT 0 248.815 0.070 248.885 ;
    RECT 0 248.955 0.070 249.025 ;
    RECT 0 249.095 0.070 249.165 ;
    RECT 0 249.235 0.070 249.305 ;
    RECT 0 249.375 0.070 249.445 ;
    RECT 0 249.515 0.070 249.585 ;
    RECT 0 249.655 0.070 249.725 ;
    RECT 0 249.795 0.070 249.865 ;
    RECT 0 249.935 0.070 250.005 ;
    RECT 0 250.075 0.070 250.145 ;
    RECT 0 250.215 0.070 250.285 ;
    RECT 0 250.355 0.070 250.425 ;
    RECT 0 250.495 0.070 250.565 ;
    RECT 0 250.635 0.070 250.705 ;
    RECT 0 250.775 0.070 250.845 ;
    RECT 0 250.915 0.070 250.985 ;
    RECT 0 251.055 0.070 251.125 ;
    RECT 0 251.195 0.070 251.265 ;
    RECT 0 251.335 0.070 251.405 ;
    RECT 0 251.475 0.070 251.545 ;
    RECT 0 251.615 0.070 251.685 ;
    RECT 0 251.755 0.070 251.825 ;
    RECT 0 251.895 0.070 251.965 ;
    RECT 0 252.035 0.070 252.105 ;
    RECT 0 252.175 0.070 252.245 ;
    RECT 0 252.315 0.070 252.385 ;
    RECT 0 252.455 0.070 252.525 ;
    RECT 0 252.595 0.070 252.665 ;
    RECT 0 252.735 0.070 252.805 ;
    RECT 0 252.875 0.070 252.945 ;
    RECT 0 253.015 0.070 253.085 ;
    RECT 0 253.155 0.070 253.225 ;
    RECT 0 253.295 0.070 253.365 ;
    RECT 0 253.435 0.070 253.505 ;
    RECT 0 253.575 0.070 253.645 ;
    RECT 0 253.715 0.070 253.785 ;
    RECT 0 253.855 0.070 253.925 ;
    RECT 0 253.995 0.070 254.065 ;
    RECT 0 254.135 0.070 254.205 ;
    RECT 0 254.275 0.070 254.345 ;
    RECT 0 254.415 0.070 254.485 ;
    RECT 0 254.555 0.070 254.625 ;
    RECT 0 254.695 0.070 254.765 ;
    RECT 0 254.835 0.070 254.905 ;
    RECT 0 254.975 0.070 255.045 ;
    RECT 0 255.115 0.070 255.185 ;
    RECT 0 255.255 0.070 255.325 ;
    RECT 0 255.395 0.070 255.465 ;
    RECT 0 255.535 0.070 255.605 ;
    RECT 0 255.675 0.070 255.745 ;
    RECT 0 255.815 0.070 255.885 ;
    RECT 0 255.955 0.070 256.025 ;
    RECT 0 256.095 0.070 256.165 ;
    RECT 0 256.235 0.070 256.305 ;
    RECT 0 256.375 0.070 256.445 ;
    RECT 0 256.515 0.070 256.585 ;
    RECT 0 256.655 0.070 256.725 ;
    RECT 0 256.795 0.070 256.865 ;
    RECT 0 256.935 0.070 257.005 ;
    RECT 0 257.075 0.070 257.145 ;
    RECT 0 257.215 0.070 257.285 ;
    RECT 0 257.355 0.070 257.425 ;
    RECT 0 257.495 0.070 257.565 ;
    RECT 0 257.635 0.070 257.705 ;
    RECT 0 257.775 0.070 257.845 ;
    RECT 0 257.915 0.070 257.985 ;
    RECT 0 258.055 0.070 258.125 ;
    RECT 0 258.195 0.070 258.265 ;
    RECT 0 258.335 0.070 258.405 ;
    RECT 0 258.475 0.070 258.545 ;
    RECT 0 258.615 0.070 258.685 ;
    RECT 0 258.755 0.070 258.825 ;
    RECT 0 258.895 0.070 258.965 ;
    RECT 0 259.035 0.070 259.105 ;
    RECT 0 259.175 0.070 259.245 ;
    RECT 0 259.315 0.070 259.385 ;
    RECT 0 259.455 0.070 259.525 ;
    RECT 0 259.595 0.070 259.665 ;
    RECT 0 259.735 0.070 259.805 ;
    RECT 0 259.875 0.070 259.945 ;
    RECT 0 260.015 0.070 260.085 ;
    RECT 0 260.155 0.070 260.225 ;
    RECT 0 260.295 0.070 260.365 ;
    RECT 0 260.435 0.070 260.505 ;
    RECT 0 260.575 0.070 260.645 ;
    RECT 0 260.715 0.070 260.785 ;
    RECT 0 260.855 0.070 260.925 ;
    RECT 0 260.995 0.070 261.065 ;
    RECT 0 261.135 0.070 261.205 ;
    RECT 0 261.275 0.070 261.345 ;
    RECT 0 261.415 0.070 261.485 ;
    RECT 0 261.555 0.070 261.625 ;
    RECT 0 261.695 0.070 261.765 ;
    RECT 0 261.835 0.070 261.905 ;
    RECT 0 261.975 0.070 262.045 ;
    RECT 0 262.115 0.070 262.185 ;
    RECT 0 262.255 0.070 262.325 ;
    RECT 0 262.395 0.070 262.465 ;
    RECT 0 262.535 0.070 262.605 ;
    RECT 0 262.675 0.070 262.745 ;
    RECT 0 262.815 0.070 262.885 ;
    RECT 0 262.955 0.070 263.025 ;
    RECT 0 263.095 0.070 263.165 ;
    RECT 0 263.235 0.070 263.305 ;
    RECT 0 263.375 0.070 263.445 ;
    RECT 0 263.515 0.070 263.585 ;
    RECT 0 263.655 0.070 263.725 ;
    RECT 0 263.795 0.070 263.865 ;
    RECT 0 263.935 0.070 264.005 ;
    RECT 0 264.075 0.070 264.145 ;
    RECT 0 264.215 0.070 264.285 ;
    RECT 0 264.355 0.070 264.425 ;
    RECT 0 264.495 0.070 264.565 ;
    RECT 0 264.635 0.070 264.705 ;
    RECT 0 264.775 0.070 264.845 ;
    RECT 0 264.915 0.070 264.985 ;
    RECT 0 265.055 0.070 265.125 ;
    RECT 0 265.195 0.070 265.265 ;
    RECT 0 265.335 0.070 265.405 ;
    RECT 0 265.475 0.070 265.545 ;
    RECT 0 265.615 0.070 265.685 ;
    RECT 0 265.755 0.070 265.825 ;
    RECT 0 265.895 0.070 265.965 ;
    RECT 0 266.035 0.070 266.105 ;
    RECT 0 266.175 0.070 266.245 ;
    RECT 0 266.315 0.070 266.385 ;
    RECT 0 266.455 0.070 266.525 ;
    RECT 0 266.595 0.070 266.665 ;
    RECT 0 266.735 0.070 266.805 ;
    RECT 0 266.875 0.070 266.945 ;
    RECT 0 267.015 0.070 267.085 ;
    RECT 0 267.155 0.070 267.225 ;
    RECT 0 267.295 0.070 267.365 ;
    RECT 0 267.435 0.070 267.505 ;
    RECT 0 267.575 0.070 267.645 ;
    RECT 0 267.715 0.070 267.785 ;
    RECT 0 267.855 0.070 267.925 ;
    RECT 0 267.995 0.070 268.065 ;
    RECT 0 268.135 0.070 268.205 ;
    RECT 0 268.275 0.070 268.345 ;
    RECT 0 268.415 0.070 268.485 ;
    RECT 0 268.555 0.070 268.625 ;
    RECT 0 268.695 0.070 268.765 ;
    RECT 0 268.835 0.070 268.905 ;
    RECT 0 268.975 0.070 269.045 ;
    RECT 0 269.115 0.070 269.185 ;
    RECT 0 269.255 0.070 269.325 ;
    RECT 0 269.395 0.070 269.465 ;
    RECT 0 269.535 0.070 269.605 ;
    RECT 0 269.675 0.070 269.745 ;
    RECT 0 269.815 0.070 269.885 ;
    RECT 0 269.955 0.070 270.025 ;
    RECT 0 270.095 0.070 270.165 ;
    RECT 0 270.235 0.070 270.305 ;
    RECT 0 270.375 0.070 270.445 ;
    RECT 0 270.515 0.070 270.585 ;
    RECT 0 270.655 0.070 270.725 ;
    RECT 0 270.795 0.070 270.865 ;
    RECT 0 270.935 0.070 271.005 ;
    RECT 0 271.075 0.070 271.145 ;
    RECT 0 271.215 0.070 271.285 ;
    RECT 0 271.355 0.070 271.425 ;
    RECT 0 271.495 0.070 271.565 ;
    RECT 0 271.635 0.070 271.705 ;
    RECT 0 271.775 0.070 271.845 ;
    RECT 0 271.915 0.070 271.985 ;
    RECT 0 272.055 0.070 272.125 ;
    RECT 0 272.195 0.070 272.265 ;
    RECT 0 272.335 0.070 272.405 ;
    RECT 0 272.475 0.070 272.545 ;
    RECT 0 272.615 0.070 272.685 ;
    RECT 0 272.755 0.070 272.825 ;
    RECT 0 272.895 0.070 272.965 ;
    RECT 0 273.035 0.070 273.105 ;
    RECT 0 273.175 0.070 273.245 ;
    RECT 0 273.315 0.070 273.385 ;
    RECT 0 273.455 0.070 273.525 ;
    RECT 0 273.595 0.070 273.665 ;
    RECT 0 273.735 0.070 273.805 ;
    RECT 0 273.875 0.070 273.945 ;
    RECT 0 274.015 0.070 274.085 ;
    RECT 0 274.155 0.070 274.225 ;
    RECT 0 274.295 0.070 274.365 ;
    RECT 0 274.435 0.070 274.505 ;
    RECT 0 274.575 0.070 274.645 ;
    RECT 0 274.715 0.070 274.785 ;
    RECT 0 274.855 0.070 274.925 ;
    RECT 0 274.995 0.070 275.065 ;
    RECT 0 275.135 0.070 275.205 ;
    RECT 0 275.275 0.070 275.345 ;
    RECT 0 275.415 0.070 275.485 ;
    RECT 0 275.555 0.070 275.625 ;
    RECT 0 275.695 0.070 275.765 ;
    RECT 0 275.835 0.070 275.905 ;
    RECT 0 275.975 0.070 276.045 ;
    RECT 0 276.115 0.070 276.185 ;
    RECT 0 276.255 0.070 276.325 ;
    RECT 0 276.395 0.070 276.465 ;
    RECT 0 276.535 0.070 276.605 ;
    RECT 0 276.675 0.070 276.745 ;
    RECT 0 276.815 0.070 276.885 ;
    RECT 0 276.955 0.070 277.025 ;
    RECT 0 277.095 0.070 277.165 ;
    RECT 0 277.235 0.070 277.305 ;
    RECT 0 277.375 0.070 277.445 ;
    RECT 0 277.515 0.070 277.585 ;
    RECT 0 277.655 0.070 277.725 ;
    RECT 0 277.795 0.070 277.865 ;
    RECT 0 277.935 0.070 278.005 ;
    RECT 0 278.075 0.070 278.145 ;
    RECT 0 278.215 0.070 278.285 ;
    RECT 0 278.355 0.070 278.425 ;
    RECT 0 278.495 0.070 278.565 ;
    RECT 0 278.635 0.070 278.705 ;
    RECT 0 278.775 0.070 278.845 ;
    RECT 0 278.915 0.070 278.985 ;
    RECT 0 279.055 0.070 279.125 ;
    RECT 0 279.195 0.070 279.265 ;
    RECT 0 279.335 0.070 279.405 ;
    RECT 0 279.475 0.070 279.545 ;
    RECT 0 279.615 0.070 279.685 ;
    RECT 0 279.755 0.070 279.825 ;
    RECT 0 279.895 0.070 279.965 ;
    RECT 0 280.035 0.070 280.105 ;
    RECT 0 280.175 0.070 280.245 ;
    RECT 0 280.315 0.070 280.385 ;
    RECT 0 280.455 0.070 280.525 ;
    RECT 0 280.595 0.070 280.665 ;
    RECT 0 280.735 0.070 280.805 ;
    RECT 0 280.875 0.070 280.945 ;
    RECT 0 281.015 0.070 281.085 ;
    RECT 0 281.155 0.070 281.225 ;
    RECT 0 281.295 0.070 281.365 ;
    RECT 0 281.435 0.070 281.505 ;
    RECT 0 281.575 0.070 281.645 ;
    RECT 0 281.715 0.070 281.785 ;
    RECT 0 281.855 0.070 281.925 ;
    RECT 0 281.995 0.070 282.065 ;
    RECT 0 282.135 0.070 282.205 ;
    RECT 0 282.275 0.070 282.345 ;
    RECT 0 282.415 0.070 282.485 ;
    RECT 0 282.555 0.070 282.625 ;
    RECT 0 282.695 0.070 282.765 ;
    RECT 0 282.835 0.070 282.905 ;
    RECT 0 282.975 0.070 283.045 ;
    RECT 0 283.115 0.070 283.185 ;
    RECT 0 283.255 0.070 283.325 ;
    RECT 0 283.395 0.070 283.465 ;
    RECT 0 283.535 0.070 283.605 ;
    RECT 0 283.675 0.070 283.745 ;
    RECT 0 283.815 0.070 283.885 ;
    RECT 0 283.955 0.070 284.025 ;
    RECT 0 284.095 0.070 284.165 ;
    RECT 0 284.235 0.070 284.305 ;
    RECT 0 284.375 0.070 284.445 ;
    RECT 0 284.515 0.070 284.585 ;
    RECT 0 284.655 0.070 284.725 ;
    RECT 0 284.795 0.070 284.865 ;
    RECT 0 284.935 0.070 285.005 ;
    RECT 0 285.075 0.070 285.145 ;
    RECT 0 285.215 0.070 285.285 ;
    RECT 0 285.355 0.070 285.425 ;
    RECT 0 285.495 0.070 285.565 ;
    RECT 0 285.635 0.070 285.705 ;
    RECT 0 285.775 0.070 285.845 ;
    RECT 0 285.915 0.070 285.985 ;
    RECT 0 286.055 0.070 286.125 ;
    RECT 0 286.195 0.070 286.265 ;
    RECT 0 286.335 0.070 286.405 ;
    RECT 0 286.475 0.070 286.545 ;
    RECT 0 286.615 0.070 286.685 ;
    RECT 0 286.755 0.070 286.825 ;
    RECT 0 286.895 0.070 286.965 ;
    RECT 0 287.035 0.070 287.105 ;
    RECT 0 287.175 0.070 287.245 ;
    RECT 0 287.315 0.070 287.385 ;
    RECT 0 287.455 0.070 287.525 ;
    RECT 0 287.595 0.070 287.665 ;
    RECT 0 287.735 0.070 287.805 ;
    RECT 0 287.875 0.070 287.945 ;
    RECT 0 288.015 0.070 288.085 ;
    RECT 0 288.155 0.070 288.225 ;
    RECT 0 288.295 0.070 288.365 ;
    RECT 0 288.435 0.070 288.505 ;
    RECT 0 288.575 0.070 288.645 ;
    RECT 0 288.715 0.070 288.785 ;
    RECT 0 288.855 0.070 288.925 ;
    RECT 0 288.995 0.070 289.065 ;
    RECT 0 289.135 0.070 289.205 ;
    RECT 0 289.275 0.070 289.345 ;
    RECT 0 289.415 0.070 289.485 ;
    RECT 0 289.555 0.070 289.625 ;
    RECT 0 289.695 0.070 289.765 ;
    RECT 0 289.835 0.070 289.905 ;
    RECT 0 289.975 0.070 290.045 ;
    RECT 0 290.115 0.070 290.185 ;
    RECT 0 290.255 0.070 290.325 ;
    RECT 0 290.395 0.070 290.465 ;
    RECT 0 290.535 0.070 290.605 ;
    RECT 0 290.675 0.070 290.745 ;
    RECT 0 290.815 0.070 290.885 ;
    RECT 0 290.955 0.070 291.025 ;
    RECT 0 291.095 0.070 291.165 ;
    RECT 0 291.235 0.070 291.305 ;
    RECT 0 291.375 0.070 291.445 ;
    RECT 0 291.515 0.070 291.585 ;
    RECT 0 291.655 0.070 291.725 ;
    RECT 0 291.795 0.070 291.865 ;
    RECT 0 291.935 0.070 292.005 ;
    RECT 0 292.075 0.070 292.145 ;
    RECT 0 292.215 0.070 292.285 ;
    RECT 0 292.355 0.070 292.425 ;
    RECT 0 292.495 0.070 292.565 ;
    RECT 0 292.635 0.070 292.705 ;
    RECT 0 292.775 0.070 292.845 ;
    RECT 0 292.915 0.070 292.985 ;
    RECT 0 293.055 0.070 293.125 ;
    RECT 0 293.195 0.070 293.265 ;
    RECT 0 293.335 0.070 293.405 ;
    RECT 0 293.475 0.070 293.545 ;
    RECT 0 293.615 0.070 293.685 ;
    RECT 0 293.755 0.070 293.825 ;
    RECT 0 293.895 0.070 293.965 ;
    RECT 0 294.035 0.070 294.105 ;
    RECT 0 294.175 0.070 294.245 ;
    RECT 0 294.315 0.070 294.385 ;
    RECT 0 294.455 0.070 294.525 ;
    RECT 0 294.595 0.070 294.665 ;
    RECT 0 294.735 0.070 294.805 ;
    RECT 0 294.875 0.070 294.945 ;
    RECT 0 295.015 0.070 295.085 ;
    RECT 0 295.155 0.070 295.225 ;
    RECT 0 295.295 0.070 295.365 ;
    RECT 0 295.435 0.070 295.505 ;
    RECT 0 295.575 0.070 295.645 ;
    RECT 0 295.715 0.070 295.785 ;
    RECT 0 295.855 0.070 295.925 ;
    RECT 0 295.995 0.070 296.065 ;
    RECT 0 296.135 0.070 296.205 ;
    RECT 0 296.275 0.070 296.345 ;
    RECT 0 296.415 0.070 296.485 ;
    RECT 0 296.555 0.070 296.625 ;
    RECT 0 296.695 0.070 296.765 ;
    RECT 0 296.835 0.070 296.905 ;
    RECT 0 296.975 0.070 297.045 ;
    RECT 0 297.115 0.070 297.185 ;
    RECT 0 297.255 0.070 297.325 ;
    RECT 0 297.395 0.070 297.465 ;
    RECT 0 297.535 0.070 297.605 ;
    RECT 0 297.675 0.070 297.745 ;
    RECT 0 297.815 0.070 297.885 ;
    RECT 0 297.955 0.070 298.025 ;
    RECT 0 298.095 0.070 298.165 ;
    RECT 0 298.235 0.070 298.305 ;
    RECT 0 298.375 0.070 298.445 ;
    RECT 0 298.515 0.070 298.585 ;
    RECT 0 298.655 0.070 298.725 ;
    RECT 0 298.795 0.070 298.865 ;
    RECT 0 298.935 0.070 299.005 ;
    RECT 0 299.075 0.070 299.145 ;
    RECT 0 299.215 0.070 299.285 ;
    RECT 0 299.355 0.070 299.425 ;
    RECT 0 299.495 0.070 299.565 ;
    RECT 0 299.635 0.070 299.705 ;
    RECT 0 299.775 0.070 299.845 ;
    RECT 0 299.915 0.070 299.985 ;
    RECT 0 300.055 0.070 300.125 ;
    RECT 0 300.195 0.070 300.265 ;
    RECT 0 300.335 0.070 300.405 ;
    RECT 0 300.475 0.070 300.545 ;
    RECT 0 300.615 0.070 300.685 ;
    RECT 0 300.755 0.070 300.825 ;
    RECT 0 300.895 0.070 300.965 ;
    RECT 0 301.035 0.070 301.105 ;
    RECT 0 301.175 0.070 301.245 ;
    RECT 0 301.315 0.070 301.385 ;
    RECT 0 301.455 0.070 301.525 ;
    RECT 0 301.595 0.070 301.665 ;
    RECT 0 301.735 0.070 301.805 ;
    RECT 0 301.875 0.070 301.945 ;
    RECT 0 302.015 0.070 302.085 ;
    RECT 0 302.155 0.070 302.225 ;
    RECT 0 302.295 0.070 302.365 ;
    RECT 0 302.435 0.070 302.505 ;
    RECT 0 302.575 0.070 302.645 ;
    RECT 0 302.715 0.070 302.785 ;
    RECT 0 302.855 0.070 302.925 ;
    RECT 0 302.995 0.070 303.065 ;
    RECT 0 303.135 0.070 303.205 ;
    RECT 0 303.275 0.070 303.345 ;
    RECT 0 303.415 0.070 303.485 ;
    RECT 0 303.555 0.070 303.625 ;
    RECT 0 303.695 0.070 303.765 ;
    RECT 0 303.835 0.070 303.905 ;
    RECT 0 303.975 0.070 304.045 ;
    RECT 0 304.115 0.070 304.185 ;
    RECT 0 304.255 0.070 304.325 ;
    RECT 0 304.395 0.070 304.465 ;
    RECT 0 304.535 0.070 304.605 ;
    RECT 0 304.675 0.070 304.745 ;
    RECT 0 304.815 0.070 304.885 ;
    RECT 0 304.955 0.070 305.025 ;
    RECT 0 305.095 0.070 305.165 ;
    RECT 0 305.235 0.070 305.305 ;
    RECT 0 305.375 0.070 305.445 ;
    RECT 0 305.515 0.070 305.585 ;
    RECT 0 305.655 0.070 305.725 ;
    RECT 0 305.795 0.070 305.865 ;
    RECT 0 305.935 0.070 306.005 ;
    RECT 0 306.075 0.070 306.145 ;
    RECT 0 306.215 0.070 306.285 ;
    RECT 0 306.355 0.070 306.425 ;
    RECT 0 306.495 0.070 306.565 ;
    RECT 0 306.635 0.070 306.705 ;
    RECT 0 306.775 0.070 306.845 ;
    RECT 0 306.915 0.070 306.985 ;
    RECT 0 307.055 0.070 307.125 ;
    RECT 0 307.195 0.070 307.265 ;
    RECT 0 307.335 0.070 307.405 ;
    RECT 0 307.475 0.070 307.545 ;
    RECT 0 307.615 0.070 307.685 ;
    RECT 0 307.755 0.070 307.825 ;
    RECT 0 307.895 0.070 307.965 ;
    RECT 0 308.035 0.070 308.105 ;
    RECT 0 308.175 0.070 308.245 ;
    RECT 0 308.315 0.070 308.385 ;
    RECT 0 308.455 0.070 308.525 ;
    RECT 0 308.595 0.070 308.665 ;
    RECT 0 308.735 0.070 308.805 ;
    RECT 0 308.875 0.070 308.945 ;
    RECT 0 309.015 0.070 309.085 ;
    RECT 0 309.155 0.070 309.225 ;
    RECT 0 309.295 0.070 309.365 ;
    RECT 0 309.435 0.070 309.505 ;
    RECT 0 309.575 0.070 309.645 ;
    RECT 0 309.715 0.070 309.785 ;
    RECT 0 309.855 0.070 309.925 ;
    RECT 0 309.995 0.070 310.065 ;
    RECT 0 310.135 0.070 310.205 ;
    RECT 0 310.275 0.070 310.345 ;
    RECT 0 310.415 0.070 310.485 ;
    RECT 0 310.555 0.070 310.625 ;
    RECT 0 310.695 0.070 310.765 ;
    RECT 0 310.835 0.070 310.905 ;
    RECT 0 310.975 0.070 311.045 ;
    RECT 0 311.115 0.070 311.185 ;
    RECT 0 311.255 0.070 311.325 ;
    RECT 0 311.395 0.070 311.465 ;
    RECT 0 311.535 0.070 311.605 ;
    RECT 0 311.675 0.070 311.745 ;
    RECT 0 311.815 0.070 311.885 ;
    RECT 0 311.955 0.070 312.025 ;
    RECT 0 312.095 0.070 312.165 ;
    RECT 0 312.235 0.070 312.305 ;
    RECT 0 312.375 0.070 312.445 ;
    RECT 0 312.515 0.070 312.585 ;
    RECT 0 312.655 0.070 312.725 ;
    RECT 0 312.795 0.070 312.865 ;
    RECT 0 312.935 0.070 313.005 ;
    RECT 0 313.075 0.070 313.145 ;
    RECT 0 313.215 0.070 313.285 ;
    RECT 0 313.355 0.070 313.425 ;
    RECT 0 313.495 0.070 313.565 ;
    RECT 0 313.635 0.070 313.705 ;
    RECT 0 313.775 0.070 313.845 ;
    RECT 0 313.915 0.070 313.985 ;
    RECT 0 314.055 0.070 314.125 ;
    RECT 0 314.195 0.070 314.265 ;
    RECT 0 314.335 0.070 314.405 ;
    RECT 0 314.475 0.070 314.545 ;
    RECT 0 314.615 0.070 314.685 ;
    RECT 0 314.755 0.070 314.825 ;
    RECT 0 314.895 0.070 314.965 ;
    RECT 0 315.035 0.070 315.105 ;
    RECT 0 315.175 0.070 315.245 ;
    RECT 0 315.315 0.070 315.385 ;
    RECT 0 315.455 0.070 315.525 ;
    RECT 0 315.595 0.070 315.665 ;
    RECT 0 315.735 0.070 315.805 ;
    RECT 0 315.875 0.070 315.945 ;
    RECT 0 316.015 0.070 316.085 ;
    RECT 0 316.155 0.070 316.225 ;
    RECT 0 316.295 0.070 316.365 ;
    RECT 0 316.435 0.070 316.505 ;
    RECT 0 316.575 0.070 316.645 ;
    RECT 0 316.715 0.070 316.785 ;
    RECT 0 316.855 0.070 316.925 ;
    RECT 0 316.995 0.070 317.065 ;
    RECT 0 317.135 0.070 317.205 ;
    RECT 0 317.275 0.070 317.345 ;
    RECT 0 317.415 0.070 317.485 ;
    RECT 0 317.555 0.070 317.625 ;
    RECT 0 317.695 0.070 317.765 ;
    RECT 0 317.835 0.070 317.905 ;
    RECT 0 317.975 0.070 318.045 ;
    RECT 0 318.115 0.070 318.185 ;
    RECT 0 318.255 0.070 318.325 ;
    RECT 0 318.395 0.070 318.465 ;
    RECT 0 318.535 0.070 318.605 ;
    RECT 0 318.675 0.070 318.745 ;
    RECT 0 318.815 0.070 318.885 ;
    RECT 0 318.955 0.070 319.025 ;
    RECT 0 319.095 0.070 319.165 ;
    RECT 0 319.235 0.070 319.305 ;
    RECT 0 319.375 0.070 319.445 ;
    RECT 0 319.515 0.070 319.585 ;
    RECT 0 319.655 0.070 319.725 ;
    RECT 0 319.795 0.070 319.865 ;
    RECT 0 319.935 0.070 320.005 ;
    RECT 0 320.075 0.070 320.145 ;
    RECT 0 320.215 0.070 320.285 ;
    RECT 0 320.355 0.070 320.425 ;
    RECT 0 320.495 0.070 320.565 ;
    RECT 0 320.635 0.070 320.705 ;
    RECT 0 320.775 0.070 320.845 ;
    RECT 0 320.915 0.070 320.985 ;
    RECT 0 321.055 0.070 321.125 ;
    RECT 0 321.195 0.070 321.265 ;
    RECT 0 321.335 0.070 321.405 ;
    RECT 0 321.475 0.070 321.545 ;
    RECT 0 321.615 0.070 321.685 ;
    RECT 0 321.755 0.070 321.825 ;
    RECT 0 321.895 0.070 321.965 ;
    RECT 0 322.035 0.070 322.105 ;
    RECT 0 322.175 0.070 322.245 ;
    RECT 0 322.315 0.070 322.385 ;
    RECT 0 322.455 0.070 322.525 ;
    RECT 0 322.595 0.070 322.665 ;
    RECT 0 322.735 0.070 322.805 ;
    RECT 0 322.875 0.070 322.945 ;
    RECT 0 323.015 0.070 323.085 ;
    RECT 0 323.155 0.070 323.225 ;
    RECT 0 323.295 0.070 323.365 ;
    RECT 0 323.435 0.070 323.505 ;
    RECT 0 323.575 0.070 323.645 ;
    RECT 0 323.715 0.070 323.785 ;
    RECT 0 323.855 0.070 323.925 ;
    RECT 0 323.995 0.070 324.065 ;
    RECT 0 324.135 0.070 324.205 ;
    RECT 0 324.275 0.070 324.345 ;
    RECT 0 324.415 0.070 324.485 ;
    RECT 0 324.555 0.070 324.625 ;
    RECT 0 324.695 0.070 324.765 ;
    RECT 0 324.835 0.070 324.905 ;
    RECT 0 324.975 0.070 325.045 ;
    RECT 0 325.115 0.070 325.185 ;
    RECT 0 325.255 0.070 325.325 ;
    RECT 0 325.395 0.070 325.465 ;
    RECT 0 325.535 0.070 325.605 ;
    RECT 0 325.675 0.070 325.745 ;
    RECT 0 325.815 0.070 325.885 ;
    RECT 0 325.955 0.070 326.025 ;
    RECT 0 326.095 0.070 326.165 ;
    RECT 0 326.235 0.070 326.305 ;
    RECT 0 326.375 0.070 326.445 ;
    RECT 0 326.515 0.070 326.585 ;
    RECT 0 326.655 0.070 326.725 ;
    RECT 0 326.795 0.070 326.865 ;
    RECT 0 326.935 0.070 327.005 ;
    RECT 0 327.075 0.070 327.145 ;
    RECT 0 327.215 0.070 327.285 ;
    RECT 0 327.355 0.070 327.425 ;
    RECT 0 327.495 0.070 327.565 ;
    RECT 0 327.635 0.070 327.705 ;
    RECT 0 327.775 0.070 327.845 ;
    RECT 0 327.915 0.070 327.985 ;
    RECT 0 328.055 0.070 328.125 ;
    RECT 0 328.195 0.070 328.265 ;
    RECT 0 328.335 0.070 328.405 ;
    RECT 0 328.475 0.070 328.545 ;
    RECT 0 328.615 0.070 328.685 ;
    RECT 0 328.755 0.070 328.825 ;
    RECT 0 328.895 0.070 328.965 ;
    RECT 0 329.035 0.070 329.105 ;
    RECT 0 329.175 0.070 329.245 ;
    RECT 0 329.315 0.070 329.385 ;
    RECT 0 329.455 0.070 329.525 ;
    RECT 0 329.595 0.070 329.665 ;
    RECT 0 329.735 0.070 329.805 ;
    RECT 0 329.875 0.070 329.945 ;
    RECT 0 330.015 0.070 330.085 ;
    RECT 0 330.155 0.070 330.225 ;
    RECT 0 330.295 0.070 330.365 ;
    RECT 0 330.435 0.070 330.505 ;
    RECT 0 330.575 0.070 330.645 ;
    RECT 0 330.715 0.070 330.785 ;
    RECT 0 330.855 0.070 330.925 ;
    RECT 0 330.995 0.070 331.065 ;
    RECT 0 331.135 0.070 331.205 ;
    RECT 0 331.275 0.070 331.345 ;
    RECT 0 331.415 0.070 331.485 ;
    RECT 0 331.555 0.070 331.625 ;
    RECT 0 331.695 0.070 331.765 ;
    RECT 0 331.835 0.070 331.905 ;
    RECT 0 331.975 0.070 332.045 ;
    RECT 0 332.115 0.070 332.185 ;
    RECT 0 332.255 0.070 332.325 ;
    RECT 0 332.395 0.070 332.465 ;
    RECT 0 332.535 0.070 332.605 ;
    RECT 0 332.675 0.070 332.745 ;
    RECT 0 332.815 0.070 332.885 ;
    RECT 0 332.955 0.070 333.025 ;
    RECT 0 333.095 0.070 333.165 ;
    RECT 0 333.235 0.070 333.305 ;
    RECT 0 333.375 0.070 333.445 ;
    RECT 0 333.515 0.070 333.585 ;
    RECT 0 333.655 0.070 333.725 ;
    RECT 0 333.795 0.070 333.865 ;
    RECT 0 333.935 0.070 334.005 ;
    RECT 0 334.075 0.070 334.145 ;
    RECT 0 334.215 0.070 334.285 ;
    RECT 0 334.355 0.070 334.425 ;
    RECT 0 334.495 0.070 334.565 ;
    RECT 0 334.635 0.070 334.705 ;
    RECT 0 334.775 0.070 334.845 ;
    RECT 0 334.915 0.070 334.985 ;
    RECT 0 335.055 0.070 335.125 ;
    RECT 0 335.195 0.070 335.265 ;
    RECT 0 335.335 0.070 335.405 ;
    RECT 0 335.475 0.070 335.545 ;
    RECT 0 335.615 0.070 335.685 ;
    RECT 0 335.755 0.070 335.825 ;
    RECT 0 335.895 0.070 335.965 ;
    RECT 0 336.035 0.070 336.105 ;
    RECT 0 336.175 0.070 336.245 ;
    RECT 0 336.315 0.070 336.385 ;
    RECT 0 336.455 0.070 336.525 ;
    RECT 0 336.595 0.070 336.665 ;
    RECT 0 336.735 0.070 336.805 ;
    RECT 0 336.875 0.070 336.945 ;
    RECT 0 337.015 0.070 337.085 ;
    RECT 0 337.155 0.070 337.225 ;
    RECT 0 337.295 0.070 337.365 ;
    RECT 0 337.435 0.070 337.505 ;
    RECT 0 337.575 0.070 337.645 ;
    RECT 0 337.715 0.070 337.785 ;
    RECT 0 337.855 0.070 337.925 ;
    RECT 0 337.995 0.070 338.065 ;
    RECT 0 338.135 0.070 338.205 ;
    RECT 0 338.275 0.070 338.345 ;
    RECT 0 338.415 0.070 338.485 ;
    RECT 0 338.555 0.070 338.625 ;
    RECT 0 338.695 0.070 338.765 ;
    RECT 0 338.835 0.070 338.905 ;
    RECT 0 338.975 0.070 339.045 ;
    RECT 0 339.115 0.070 339.185 ;
    RECT 0 339.255 0.070 339.325 ;
    RECT 0 339.395 0.070 339.465 ;
    RECT 0 339.535 0.070 339.605 ;
    RECT 0 339.675 0.070 339.745 ;
    RECT 0 339.815 0.070 339.885 ;
    RECT 0 339.955 0.070 340.025 ;
    RECT 0 340.095 0.070 340.165 ;
    RECT 0 340.235 0.070 340.305 ;
    RECT 0 340.375 0.070 340.445 ;
    RECT 0 340.515 0.070 340.585 ;
    RECT 0 340.655 0.070 340.725 ;
    RECT 0 340.795 0.070 340.865 ;
    RECT 0 340.935 0.070 341.005 ;
    RECT 0 341.075 0.070 341.145 ;
    RECT 0 341.215 0.070 341.285 ;
    RECT 0 341.355 0.070 341.425 ;
    RECT 0 341.495 0.070 341.565 ;
    RECT 0 341.635 0.070 341.705 ;
    RECT 0 341.775 0.070 341.845 ;
    RECT 0 341.915 0.070 341.985 ;
    RECT 0 342.055 0.070 342.125 ;
    RECT 0 342.195 0.070 342.265 ;
    RECT 0 342.335 0.070 342.405 ;
    RECT 0 342.475 0.070 342.545 ;
    RECT 0 342.615 0.070 342.685 ;
    RECT 0 342.755 0.070 342.825 ;
    RECT 0 342.895 0.070 342.965 ;
    RECT 0 343.035 0.070 343.105 ;
    RECT 0 343.175 0.070 343.245 ;
    RECT 0 343.315 0.070 343.385 ;
    RECT 0 343.455 0.070 343.525 ;
    RECT 0 343.595 0.070 343.665 ;
    RECT 0 343.735 0.070 343.805 ;
    RECT 0 343.875 0.070 343.945 ;
    RECT 0 344.015 0.070 344.085 ;
    RECT 0 344.155 0.070 344.225 ;
    RECT 0 344.295 0.070 344.365 ;
    RECT 0 344.435 0.070 344.505 ;
    RECT 0 344.575 0.070 344.645 ;
    RECT 0 344.715 0.070 344.785 ;
    RECT 0 344.855 0.070 344.925 ;
    RECT 0 344.995 0.070 345.065 ;
    RECT 0 345.135 0.070 345.205 ;
    RECT 0 345.275 0.070 345.345 ;
    RECT 0 345.415 0.070 345.485 ;
    RECT 0 345.555 0.070 345.625 ;
    RECT 0 345.695 0.070 345.765 ;
    RECT 0 345.835 0.070 345.905 ;
    RECT 0 345.975 0.070 346.045 ;
    RECT 0 346.115 0.070 346.185 ;
    RECT 0 346.255 0.070 346.325 ;
    RECT 0 346.395 0.070 346.465 ;
    RECT 0 346.535 0.070 346.605 ;
    RECT 0 346.675 0.070 346.745 ;
    RECT 0 346.815 0.070 346.885 ;
    RECT 0 346.955 0.070 347.025 ;
    RECT 0 347.095 0.070 347.165 ;
    RECT 0 347.235 0.070 347.305 ;
    RECT 0 347.375 0.070 347.445 ;
    RECT 0 347.515 0.070 347.585 ;
    RECT 0 347.655 0.070 347.725 ;
    RECT 0 347.795 0.070 347.865 ;
    RECT 0 347.935 0.070 348.005 ;
    RECT 0 348.075 0.070 348.145 ;
    RECT 0 348.215 0.070 348.285 ;
    RECT 0 348.355 0.070 348.425 ;
    RECT 0 348.495 0.070 348.565 ;
    RECT 0 348.635 0.070 348.705 ;
    RECT 0 348.775 0.070 348.845 ;
    RECT 0 348.915 0.070 348.985 ;
    RECT 0 349.055 0.070 349.125 ;
    RECT 0 349.195 0.070 349.265 ;
    RECT 0 349.335 0.070 349.405 ;
    RECT 0 349.475 0.070 349.545 ;
    RECT 0 349.615 0.070 349.685 ;
    RECT 0 349.755 0.070 349.825 ;
    RECT 0 349.895 0.070 349.965 ;
    RECT 0 350.035 0.070 350.105 ;
    RECT 0 350.175 0.070 350.245 ;
    RECT 0 350.315 0.070 350.385 ;
    RECT 0 350.455 0.070 350.525 ;
    RECT 0 350.595 0.070 350.665 ;
    RECT 0 350.735 0.070 350.805 ;
    RECT 0 350.875 0.070 350.945 ;
    RECT 0 351.015 0.070 351.085 ;
    RECT 0 351.155 0.070 351.225 ;
    RECT 0 351.295 0.070 351.365 ;
    RECT 0 351.435 0.070 351.505 ;
    RECT 0 351.575 0.070 351.645 ;
    RECT 0 351.715 0.070 351.785 ;
    RECT 0 351.855 0.070 351.925 ;
    RECT 0 351.995 0.070 352.065 ;
    RECT 0 352.135 0.070 352.205 ;
    RECT 0 352.275 0.070 352.345 ;
    RECT 0 352.415 0.070 352.485 ;
    RECT 0 352.555 0.070 352.625 ;
    RECT 0 352.695 0.070 352.765 ;
    RECT 0 352.835 0.070 352.905 ;
    RECT 0 352.975 0.070 353.045 ;
    RECT 0 353.115 0.070 353.185 ;
    RECT 0 353.255 0.070 353.325 ;
    RECT 0 353.395 0.070 353.465 ;
    RECT 0 353.535 0.070 353.605 ;
    RECT 0 353.675 0.070 353.745 ;
    RECT 0 353.815 0.070 353.885 ;
    RECT 0 353.955 0.070 354.025 ;
    RECT 0 354.095 0.070 354.165 ;
    RECT 0 354.235 0.070 354.305 ;
    RECT 0 354.375 0.070 354.445 ;
    RECT 0 354.515 0.070 354.585 ;
    RECT 0 354.655 0.070 354.725 ;
    RECT 0 354.795 0.070 354.865 ;
    RECT 0 354.935 0.070 355.005 ;
    RECT 0 355.075 0.070 355.145 ;
    RECT 0 355.215 0.070 355.285 ;
    RECT 0 355.355 0.070 355.425 ;
    RECT 0 355.495 0.070 355.565 ;
    RECT 0 355.635 0.070 355.705 ;
    RECT 0 355.775 0.070 355.845 ;
    RECT 0 355.915 0.070 355.985 ;
    RECT 0 356.055 0.070 356.125 ;
    RECT 0 356.195 0.070 356.265 ;
    RECT 0 356.335 0.070 356.405 ;
    RECT 0 356.475 0.070 356.545 ;
    RECT 0 356.615 0.070 356.685 ;
    RECT 0 356.755 0.070 356.825 ;
    RECT 0 356.895 0.070 356.965 ;
    RECT 0 357.035 0.070 357.105 ;
    RECT 0 357.175 0.070 357.245 ;
    RECT 0 357.315 0.070 357.385 ;
    RECT 0 357.455 0.070 357.525 ;
    RECT 0 357.595 0.070 357.665 ;
    RECT 0 357.735 0.070 357.805 ;
    RECT 0 357.875 0.070 357.945 ;
    RECT 0 358.015 0.070 358.085 ;
    RECT 0 358.155 0.070 358.225 ;
    RECT 0 358.295 0.070 358.365 ;
    RECT 0 358.435 0.070 358.505 ;
    RECT 0 358.575 0.070 358.645 ;
    RECT 0 358.715 0.070 358.785 ;
    RECT 0 358.855 0.070 358.925 ;
    RECT 0 358.995 0.070 359.065 ;
    RECT 0 359.135 0.070 359.205 ;
    RECT 0 359.275 0.070 359.345 ;
    RECT 0 359.415 0.070 359.485 ;
    RECT 0 359.555 0.070 359.625 ;
    RECT 0 359.695 0.070 359.765 ;
    RECT 0 359.835 0.070 359.905 ;
    RECT 0 359.975 0.070 360.045 ;
    RECT 0 360.115 0.070 360.185 ;
    RECT 0 360.255 0.070 360.325 ;
    RECT 0 360.395 0.070 360.465 ;
    RECT 0 360.535 0.070 360.605 ;
    RECT 0 360.675 0.070 360.745 ;
    RECT 0 360.815 0.070 360.885 ;
    RECT 0 360.955 0.070 361.025 ;
    RECT 0 361.095 0.070 361.165 ;
    RECT 0 361.235 0.070 361.305 ;
    RECT 0 361.375 0.070 361.445 ;
    RECT 0 361.515 0.070 361.585 ;
    RECT 0 361.655 0.070 361.725 ;
    RECT 0 361.795 0.070 361.865 ;
    RECT 0 361.935 0.070 362.005 ;
    RECT 0 362.075 0.070 362.145 ;
    RECT 0 362.215 0.070 362.285 ;
    RECT 0 362.355 0.070 362.425 ;
    RECT 0 362.495 0.070 362.565 ;
    RECT 0 362.635 0.070 362.705 ;
    RECT 0 362.775 0.070 362.845 ;
    RECT 0 362.915 0.070 362.985 ;
    RECT 0 363.055 0.070 363.125 ;
    RECT 0 363.195 0.070 363.265 ;
    RECT 0 363.335 0.070 363.405 ;
    RECT 0 363.475 0.070 363.545 ;
    RECT 0 363.615 0.070 363.685 ;
    RECT 0 363.755 0.070 363.825 ;
    RECT 0 363.895 0.070 363.965 ;
    RECT 0 364.035 0.070 364.105 ;
    RECT 0 364.175 0.070 364.245 ;
    RECT 0 364.315 0.070 364.385 ;
    RECT 0 364.455 0.070 364.525 ;
    RECT 0 364.595 0.070 364.665 ;
    RECT 0 364.735 0.070 364.805 ;
    RECT 0 364.875 0.070 364.945 ;
    RECT 0 365.015 0.070 365.085 ;
    RECT 0 365.155 0.070 365.225 ;
    RECT 0 365.295 0.070 365.365 ;
    RECT 0 365.435 0.070 365.505 ;
    RECT 0 365.575 0.070 365.645 ;
    RECT 0 365.715 0.070 365.785 ;
    RECT 0 365.855 0.070 365.925 ;
    RECT 0 365.995 0.070 366.065 ;
    RECT 0 366.135 0.070 366.205 ;
    RECT 0 366.275 0.070 366.345 ;
    RECT 0 366.415 0.070 366.485 ;
    RECT 0 366.555 0.070 366.625 ;
    RECT 0 366.695 0.070 366.765 ;
    RECT 0 366.835 0.070 366.905 ;
    RECT 0 366.975 0.070 367.045 ;
    RECT 0 367.115 0.070 367.185 ;
    RECT 0 367.255 0.070 367.325 ;
    RECT 0 367.395 0.070 367.465 ;
    RECT 0 367.535 0.070 367.605 ;
    RECT 0 367.675 0.070 367.745 ;
    RECT 0 367.815 0.070 367.885 ;
    RECT 0 367.955 0.070 368.025 ;
    RECT 0 368.095 0.070 368.165 ;
    RECT 0 368.235 0.070 368.305 ;
    RECT 0 368.375 0.070 368.445 ;
    RECT 0 368.515 0.070 368.585 ;
    RECT 0 368.655 0.070 368.725 ;
    RECT 0 368.795 0.070 368.865 ;
    RECT 0 368.935 0.070 369.005 ;
    RECT 0 369.075 0.070 369.145 ;
    RECT 0 369.215 0.070 369.285 ;
    RECT 0 369.355 0.070 369.425 ;
    RECT 0 369.495 0.070 369.565 ;
    RECT 0 369.635 0.070 369.705 ;
    RECT 0 369.775 0.070 369.845 ;
    RECT 0 369.915 0.070 369.985 ;
    RECT 0 370.055 0.070 370.125 ;
    RECT 0 370.195 0.070 370.265 ;
    RECT 0 370.335 0.070 370.405 ;
    RECT 0 370.475 0.070 370.545 ;
    RECT 0 370.615 0.070 370.685 ;
    RECT 0 370.755 0.070 370.825 ;
    RECT 0 370.895 0.070 370.965 ;
    RECT 0 371.035 0.070 371.105 ;
    RECT 0 371.175 0.070 371.245 ;
    RECT 0 371.315 0.070 371.385 ;
    RECT 0 371.455 0.070 371.525 ;
    RECT 0 371.595 0.070 371.665 ;
    RECT 0 371.735 0.070 371.805 ;
    RECT 0 371.875 0.070 371.945 ;
    RECT 0 372.015 0.070 372.085 ;
    RECT 0 372.155 0.070 372.225 ;
    RECT 0 372.295 0.070 372.365 ;
    RECT 0 372.435 0.070 372.505 ;
    RECT 0 372.575 0.070 372.645 ;
    RECT 0 372.715 0.070 372.785 ;
    RECT 0 372.855 0.070 372.925 ;
    RECT 0 372.995 0.070 373.065 ;
    RECT 0 373.135 0.070 373.205 ;
    RECT 0 373.275 0.070 373.345 ;
    RECT 0 373.415 0.070 373.485 ;
    RECT 0 373.555 0.070 373.625 ;
    RECT 0 373.695 0.070 373.765 ;
    RECT 0 373.835 0.070 373.905 ;
    RECT 0 373.975 0.070 374.045 ;
    RECT 0 374.115 0.070 374.185 ;
    RECT 0 374.255 0.070 374.325 ;
    RECT 0 374.395 0.070 374.465 ;
    RECT 0 374.535 0.070 374.605 ;
    RECT 0 374.675 0.070 374.745 ;
    RECT 0 374.815 0.070 374.885 ;
    RECT 0 374.955 0.070 375.025 ;
    RECT 0 375.095 0.070 375.165 ;
    RECT 0 375.235 0.070 375.305 ;
    RECT 0 375.375 0.070 375.445 ;
    RECT 0 375.515 0.070 375.585 ;
    RECT 0 375.655 0.070 375.725 ;
    RECT 0 375.795 0.070 375.865 ;
    RECT 0 375.935 0.070 376.005 ;
    RECT 0 376.075 0.070 376.145 ;
    RECT 0 376.215 0.070 376.285 ;
    RECT 0 376.355 0.070 376.425 ;
    RECT 0 376.495 0.070 376.565 ;
    RECT 0 376.635 0.070 376.705 ;
    RECT 0 376.775 0.070 376.845 ;
    RECT 0 376.915 0.070 376.985 ;
    RECT 0 377.055 0.070 377.125 ;
    RECT 0 377.195 0.070 377.265 ;
    RECT 0 377.335 0.070 377.405 ;
    RECT 0 377.475 0.070 377.545 ;
    RECT 0 377.615 0.070 377.685 ;
    RECT 0 377.755 0.070 377.825 ;
    RECT 0 377.895 0.070 377.965 ;
    RECT 0 378.035 0.070 378.105 ;
    RECT 0 378.175 0.070 378.245 ;
    RECT 0 378.315 0.070 378.385 ;
    RECT 0 378.455 0.070 378.525 ;
    RECT 0 378.595 0.070 378.665 ;
    RECT 0 378.735 0.070 378.805 ;
    RECT 0 378.875 0.070 378.945 ;
    RECT 0 379.015 0.070 379.085 ;
    RECT 0 379.155 0.070 379.225 ;
    RECT 0 379.295 0.070 379.365 ;
    RECT 0 379.435 0.070 379.505 ;
    RECT 0 379.575 0.070 379.645 ;
    RECT 0 379.715 0.070 379.785 ;
    RECT 0 379.855 0.070 379.925 ;
    RECT 0 379.995 0.070 380.065 ;
    RECT 0 380.135 0.070 380.205 ;
    RECT 0 380.275 0.070 380.345 ;
    RECT 0 380.415 0.070 380.485 ;
    RECT 0 380.555 0.070 380.625 ;
    RECT 0 380.695 0.070 380.765 ;
    RECT 0 380.835 0.070 380.905 ;
    RECT 0 380.975 0.070 381.045 ;
    RECT 0 381.115 0.070 381.185 ;
    RECT 0 381.255 0.070 381.325 ;
    RECT 0 381.395 0.070 381.465 ;
    RECT 0 381.535 0.070 381.605 ;
    RECT 0 381.675 0.070 381.745 ;
    RECT 0 381.815 0.070 381.885 ;
    RECT 0 381.955 0.070 382.025 ;
    RECT 0 382.095 0.070 382.165 ;
    RECT 0 382.235 0.070 382.305 ;
    RECT 0 382.375 0.070 382.445 ;
    RECT 0 382.515 0.070 382.585 ;
    RECT 0 382.655 0.070 382.725 ;
    RECT 0 382.795 0.070 382.865 ;
    RECT 0 382.935 0.070 383.005 ;
    RECT 0 383.075 0.070 383.145 ;
    RECT 0 383.215 0.070 383.285 ;
    RECT 0 383.355 0.070 383.425 ;
    RECT 0 383.495 0.070 383.565 ;
    RECT 0 383.635 0.070 383.705 ;
    RECT 0 383.775 0.070 383.845 ;
    RECT 0 383.915 0.070 383.985 ;
    RECT 0 384.055 0.070 384.125 ;
    RECT 0 384.195 0.070 384.265 ;
    RECT 0 384.335 0.070 384.405 ;
    RECT 0 384.475 0.070 384.545 ;
    RECT 0 384.615 0.070 384.685 ;
    RECT 0 384.755 0.070 384.825 ;
    RECT 0 384.895 0.070 384.965 ;
    RECT 0 385.035 0.070 385.105 ;
    RECT 0 385.175 0.070 385.245 ;
    RECT 0 385.315 0.070 385.385 ;
    RECT 0 385.455 0.070 385.525 ;
    RECT 0 385.595 0.070 385.665 ;
    RECT 0 385.735 0.070 385.805 ;
    RECT 0 385.875 0.070 385.945 ;
    RECT 0 386.015 0.070 386.085 ;
    RECT 0 386.155 0.070 386.225 ;
    RECT 0 386.295 0.070 386.365 ;
    RECT 0 386.435 0.070 386.505 ;
    RECT 0 386.575 0.070 386.645 ;
    RECT 0 386.715 0.070 386.785 ;
    RECT 0 386.855 0.070 386.925 ;
    RECT 0 386.995 0.070 387.065 ;
    RECT 0 387.135 0.070 387.205 ;
    RECT 0 387.275 0.070 387.345 ;
    RECT 0 387.415 0.070 387.485 ;
    RECT 0 387.555 0.070 387.625 ;
    RECT 0 387.695 0.070 387.765 ;
    RECT 0 387.835 0.070 387.905 ;
    RECT 0 387.975 0.070 388.045 ;
    RECT 0 388.115 0.070 388.185 ;
    RECT 0 388.255 0.070 388.325 ;
    RECT 0 388.395 0.070 388.465 ;
    RECT 0 388.535 0.070 388.605 ;
    RECT 0 388.675 0.070 388.745 ;
    RECT 0 388.815 0.070 388.885 ;
    RECT 0 388.955 0.070 389.025 ;
    RECT 0 389.095 0.070 389.165 ;
    RECT 0 389.235 0.070 389.305 ;
    RECT 0 389.375 0.070 389.445 ;
    RECT 0 389.515 0.070 389.585 ;
    RECT 0 389.655 0.070 389.725 ;
    RECT 0 389.795 0.070 389.865 ;
    RECT 0 389.935 0.070 390.005 ;
    RECT 0 390.075 0.070 390.145 ;
    RECT 0 390.215 0.070 390.285 ;
    RECT 0 390.355 0.070 390.425 ;
    RECT 0 390.495 0.070 390.565 ;
    RECT 0 390.635 0.070 390.705 ;
    RECT 0 390.775 0.070 390.845 ;
    RECT 0 390.915 0.070 390.985 ;
    RECT 0 391.055 0.070 391.125 ;
    RECT 0 391.195 0.070 391.265 ;
    RECT 0 391.335 0.070 391.405 ;
    RECT 0 391.475 0.070 391.545 ;
    RECT 0 391.615 0.070 391.685 ;
    RECT 0 391.755 0.070 391.825 ;
    RECT 0 391.895 0.070 391.965 ;
    RECT 0 392.035 0.070 392.105 ;
    RECT 0 392.175 0.070 392.245 ;
    RECT 0 392.315 0.070 392.385 ;
    RECT 0 392.455 0.070 392.525 ;
    RECT 0 392.595 0.070 392.665 ;
    RECT 0 392.735 0.070 392.805 ;
    RECT 0 392.875 0.070 392.945 ;
    RECT 0 393.015 0.070 393.085 ;
    RECT 0 393.155 0.070 393.225 ;
    RECT 0 393.295 0.070 393.365 ;
    RECT 0 393.435 0.070 393.505 ;
    RECT 0 393.575 0.070 393.645 ;
    RECT 0 393.715 0.070 393.785 ;
    RECT 0 393.855 0.070 393.925 ;
    RECT 0 393.995 0.070 394.065 ;
    RECT 0 394.135 0.070 394.205 ;
    RECT 0 394.275 0.070 394.345 ;
    RECT 0 394.415 0.070 394.485 ;
    RECT 0 394.555 0.070 394.625 ;
    RECT 0 394.695 0.070 394.765 ;
    RECT 0 394.835 0.070 394.905 ;
    RECT 0 394.975 0.070 395.045 ;
    RECT 0 395.115 0.070 395.185 ;
    RECT 0 395.255 0.070 395.325 ;
    RECT 0 395.395 0.070 395.465 ;
    RECT 0 395.535 0.070 395.605 ;
    RECT 0 395.675 0.070 395.745 ;
    RECT 0 395.815 0.070 395.885 ;
    RECT 0 395.955 0.070 396.025 ;
    RECT 0 396.095 0.070 396.165 ;
    RECT 0 396.235 0.070 396.305 ;
    RECT 0 396.375 0.070 396.445 ;
    RECT 0 396.515 0.070 396.585 ;
    RECT 0 396.655 0.070 396.725 ;
    RECT 0 396.795 0.070 396.865 ;
    RECT 0 396.935 0.070 397.005 ;
    RECT 0 397.075 0.070 397.145 ;
    RECT 0 397.215 0.070 397.285 ;
    RECT 0 397.355 0.070 397.425 ;
    RECT 0 397.495 0.070 397.565 ;
    RECT 0 397.635 0.070 397.705 ;
    RECT 0 397.775 0.070 397.845 ;
    RECT 0 397.915 0.070 397.985 ;
    RECT 0 398.055 0.070 398.125 ;
    RECT 0 398.195 0.070 398.265 ;
    RECT 0 398.335 0.070 398.405 ;
    RECT 0 398.475 0.070 398.545 ;
    RECT 0 398.615 0.070 398.685 ;
    RECT 0 398.755 0.070 398.825 ;
    RECT 0 398.895 0.070 398.965 ;
    RECT 0 399.035 0.070 399.105 ;
    RECT 0 399.175 0.070 399.245 ;
    RECT 0 399.315 0.070 399.385 ;
    RECT 0 399.455 0.070 399.525 ;
    RECT 0 399.595 0.070 399.665 ;
    RECT 0 399.735 0.070 399.805 ;
    RECT 0 399.875 0.070 399.945 ;
    RECT 0 400.015 0.070 504.525 ;
    RECT 0 504.595 0.070 504.665 ;
    RECT 0 504.735 0.070 504.805 ;
    RECT 0 504.875 0.070 504.945 ;
    RECT 0 505.015 0.070 505.085 ;
    RECT 0 505.155 0.070 505.225 ;
    RECT 0 505.295 0.070 505.365 ;
    RECT 0 505.435 0.070 505.505 ;
    RECT 0 505.575 0.070 505.645 ;
    RECT 0 505.715 0.070 505.785 ;
    RECT 0 505.855 0.070 505.925 ;
    RECT 0 505.995 0.070 506.065 ;
    RECT 0 506.135 0.070 506.205 ;
    RECT 0 506.275 0.070 506.345 ;
    RECT 0 506.415 0.070 506.485 ;
    RECT 0 506.555 0.070 506.625 ;
    RECT 0 506.695 0.070 506.765 ;
    RECT 0 506.835 0.070 506.905 ;
    RECT 0 506.975 0.070 507.045 ;
    RECT 0 507.115 0.070 507.185 ;
    RECT 0 507.255 0.070 507.325 ;
    RECT 0 507.395 0.070 507.465 ;
    RECT 0 507.535 0.070 507.605 ;
    RECT 0 507.675 0.070 507.745 ;
    RECT 0 507.815 0.070 507.885 ;
    RECT 0 507.955 0.070 508.025 ;
    RECT 0 508.095 0.070 508.165 ;
    RECT 0 508.235 0.070 508.305 ;
    RECT 0 508.375 0.070 508.445 ;
    RECT 0 508.515 0.070 508.585 ;
    RECT 0 508.655 0.070 508.725 ;
    RECT 0 508.795 0.070 508.865 ;
    RECT 0 508.935 0.070 509.005 ;
    RECT 0 509.075 0.070 509.145 ;
    RECT 0 509.215 0.070 509.285 ;
    RECT 0 509.355 0.070 509.425 ;
    RECT 0 509.495 0.070 509.565 ;
    RECT 0 509.635 0.070 509.705 ;
    RECT 0 509.775 0.070 509.845 ;
    RECT 0 509.915 0.070 509.985 ;
    RECT 0 510.055 0.070 510.125 ;
    RECT 0 510.195 0.070 510.265 ;
    RECT 0 510.335 0.070 510.405 ;
    RECT 0 510.475 0.070 510.545 ;
    RECT 0 510.615 0.070 510.685 ;
    RECT 0 510.755 0.070 510.825 ;
    RECT 0 510.895 0.070 510.965 ;
    RECT 0 511.035 0.070 511.105 ;
    RECT 0 511.175 0.070 511.245 ;
    RECT 0 511.315 0.070 511.385 ;
    RECT 0 511.455 0.070 511.525 ;
    RECT 0 511.595 0.070 511.665 ;
    RECT 0 511.735 0.070 511.805 ;
    RECT 0 511.875 0.070 511.945 ;
    RECT 0 512.015 0.070 512.085 ;
    RECT 0 512.155 0.070 512.225 ;
    RECT 0 512.295 0.070 512.365 ;
    RECT 0 512.435 0.070 512.505 ;
    RECT 0 512.575 0.070 512.645 ;
    RECT 0 512.715 0.070 512.785 ;
    RECT 0 512.855 0.070 512.925 ;
    RECT 0 512.995 0.070 513.065 ;
    RECT 0 513.135 0.070 513.205 ;
    RECT 0 513.275 0.070 513.345 ;
    RECT 0 513.415 0.070 513.485 ;
    RECT 0 513.555 0.070 513.625 ;
    RECT 0 513.695 0.070 513.765 ;
    RECT 0 513.835 0.070 513.905 ;
    RECT 0 513.975 0.070 514.045 ;
    RECT 0 514.115 0.070 514.185 ;
    RECT 0 514.255 0.070 514.325 ;
    RECT 0 514.395 0.070 514.465 ;
    RECT 0 514.535 0.070 514.605 ;
    RECT 0 514.675 0.070 514.745 ;
    RECT 0 514.815 0.070 514.885 ;
    RECT 0 514.955 0.070 515.025 ;
    RECT 0 515.095 0.070 515.165 ;
    RECT 0 515.235 0.070 515.305 ;
    RECT 0 515.375 0.070 515.445 ;
    RECT 0 515.515 0.070 515.585 ;
    RECT 0 515.655 0.070 515.725 ;
    RECT 0 515.795 0.070 515.865 ;
    RECT 0 515.935 0.070 516.005 ;
    RECT 0 516.075 0.070 516.145 ;
    RECT 0 516.215 0.070 516.285 ;
    RECT 0 516.355 0.070 516.425 ;
    RECT 0 516.495 0.070 516.565 ;
    RECT 0 516.635 0.070 516.705 ;
    RECT 0 516.775 0.070 516.845 ;
    RECT 0 516.915 0.070 516.985 ;
    RECT 0 517.055 0.070 517.125 ;
    RECT 0 517.195 0.070 517.265 ;
    RECT 0 517.335 0.070 517.405 ;
    RECT 0 517.475 0.070 517.545 ;
    RECT 0 517.615 0.070 517.685 ;
    RECT 0 517.755 0.070 517.825 ;
    RECT 0 517.895 0.070 517.965 ;
    RECT 0 518.035 0.070 518.105 ;
    RECT 0 518.175 0.070 518.245 ;
    RECT 0 518.315 0.070 518.385 ;
    RECT 0 518.455 0.070 518.525 ;
    RECT 0 518.595 0.070 518.665 ;
    RECT 0 518.735 0.070 518.805 ;
    RECT 0 518.875 0.070 518.945 ;
    RECT 0 519.015 0.070 519.085 ;
    RECT 0 519.155 0.070 519.225 ;
    RECT 0 519.295 0.070 519.365 ;
    RECT 0 519.435 0.070 519.505 ;
    RECT 0 519.575 0.070 519.645 ;
    RECT 0 519.715 0.070 519.785 ;
    RECT 0 519.855 0.070 519.925 ;
    RECT 0 519.995 0.070 520.065 ;
    RECT 0 520.135 0.070 520.205 ;
    RECT 0 520.275 0.070 520.345 ;
    RECT 0 520.415 0.070 520.485 ;
    RECT 0 520.555 0.070 520.625 ;
    RECT 0 520.695 0.070 520.765 ;
    RECT 0 520.835 0.070 520.905 ;
    RECT 0 520.975 0.070 521.045 ;
    RECT 0 521.115 0.070 521.185 ;
    RECT 0 521.255 0.070 521.325 ;
    RECT 0 521.395 0.070 521.465 ;
    RECT 0 521.535 0.070 521.605 ;
    RECT 0 521.675 0.070 521.745 ;
    RECT 0 521.815 0.070 521.885 ;
    RECT 0 521.955 0.070 522.025 ;
    RECT 0 522.095 0.070 522.165 ;
    RECT 0 522.235 0.070 522.305 ;
    RECT 0 522.375 0.070 522.445 ;
    RECT 0 522.515 0.070 522.585 ;
    RECT 0 522.655 0.070 522.725 ;
    RECT 0 522.795 0.070 522.865 ;
    RECT 0 522.935 0.070 523.005 ;
    RECT 0 523.075 0.070 523.145 ;
    RECT 0 523.215 0.070 523.285 ;
    RECT 0 523.355 0.070 523.425 ;
    RECT 0 523.495 0.070 523.565 ;
    RECT 0 523.635 0.070 523.705 ;
    RECT 0 523.775 0.070 523.845 ;
    RECT 0 523.915 0.070 523.985 ;
    RECT 0 524.055 0.070 524.125 ;
    RECT 0 524.195 0.070 524.265 ;
    RECT 0 524.335 0.070 524.405 ;
    RECT 0 524.475 0.070 524.545 ;
    RECT 0 524.615 0.070 524.685 ;
    RECT 0 524.755 0.070 524.825 ;
    RECT 0 524.895 0.070 524.965 ;
    RECT 0 525.035 0.070 525.105 ;
    RECT 0 525.175 0.070 525.245 ;
    RECT 0 525.315 0.070 525.385 ;
    RECT 0 525.455 0.070 525.525 ;
    RECT 0 525.595 0.070 525.665 ;
    RECT 0 525.735 0.070 525.805 ;
    RECT 0 525.875 0.070 525.945 ;
    RECT 0 526.015 0.070 526.085 ;
    RECT 0 526.155 0.070 526.225 ;
    RECT 0 526.295 0.070 526.365 ;
    RECT 0 526.435 0.070 526.505 ;
    RECT 0 526.575 0.070 526.645 ;
    RECT 0 526.715 0.070 526.785 ;
    RECT 0 526.855 0.070 526.925 ;
    RECT 0 526.995 0.070 527.065 ;
    RECT 0 527.135 0.070 527.205 ;
    RECT 0 527.275 0.070 527.345 ;
    RECT 0 527.415 0.070 527.485 ;
    RECT 0 527.555 0.070 527.625 ;
    RECT 0 527.695 0.070 527.765 ;
    RECT 0 527.835 0.070 527.905 ;
    RECT 0 527.975 0.070 528.045 ;
    RECT 0 528.115 0.070 528.185 ;
    RECT 0 528.255 0.070 528.325 ;
    RECT 0 528.395 0.070 528.465 ;
    RECT 0 528.535 0.070 528.605 ;
    RECT 0 528.675 0.070 528.745 ;
    RECT 0 528.815 0.070 528.885 ;
    RECT 0 528.955 0.070 529.025 ;
    RECT 0 529.095 0.070 529.165 ;
    RECT 0 529.235 0.070 529.305 ;
    RECT 0 529.375 0.070 529.445 ;
    RECT 0 529.515 0.070 529.585 ;
    RECT 0 529.655 0.070 529.725 ;
    RECT 0 529.795 0.070 529.865 ;
    RECT 0 529.935 0.070 530.005 ;
    RECT 0 530.075 0.070 530.145 ;
    RECT 0 530.215 0.070 530.285 ;
    RECT 0 530.355 0.070 530.425 ;
    RECT 0 530.495 0.070 530.565 ;
    RECT 0 530.635 0.070 530.705 ;
    RECT 0 530.775 0.070 530.845 ;
    RECT 0 530.915 0.070 530.985 ;
    RECT 0 531.055 0.070 531.125 ;
    RECT 0 531.195 0.070 531.265 ;
    RECT 0 531.335 0.070 531.405 ;
    RECT 0 531.475 0.070 531.545 ;
    RECT 0 531.615 0.070 531.685 ;
    RECT 0 531.755 0.070 531.825 ;
    RECT 0 531.895 0.070 531.965 ;
    RECT 0 532.035 0.070 532.105 ;
    RECT 0 532.175 0.070 532.245 ;
    RECT 0 532.315 0.070 532.385 ;
    RECT 0 532.455 0.070 532.525 ;
    RECT 0 532.595 0.070 532.665 ;
    RECT 0 532.735 0.070 532.805 ;
    RECT 0 532.875 0.070 532.945 ;
    RECT 0 533.015 0.070 533.085 ;
    RECT 0 533.155 0.070 533.225 ;
    RECT 0 533.295 0.070 533.365 ;
    RECT 0 533.435 0.070 533.505 ;
    RECT 0 533.575 0.070 533.645 ;
    RECT 0 533.715 0.070 533.785 ;
    RECT 0 533.855 0.070 533.925 ;
    RECT 0 533.995 0.070 534.065 ;
    RECT 0 534.135 0.070 534.205 ;
    RECT 0 534.275 0.070 534.345 ;
    RECT 0 534.415 0.070 534.485 ;
    RECT 0 534.555 0.070 534.625 ;
    RECT 0 534.695 0.070 534.765 ;
    RECT 0 534.835 0.070 534.905 ;
    RECT 0 534.975 0.070 535.045 ;
    RECT 0 535.115 0.070 535.185 ;
    RECT 0 535.255 0.070 535.325 ;
    RECT 0 535.395 0.070 535.465 ;
    RECT 0 535.535 0.070 535.605 ;
    RECT 0 535.675 0.070 535.745 ;
    RECT 0 535.815 0.070 535.885 ;
    RECT 0 535.955 0.070 536.025 ;
    RECT 0 536.095 0.070 536.165 ;
    RECT 0 536.235 0.070 536.305 ;
    RECT 0 536.375 0.070 536.445 ;
    RECT 0 536.515 0.070 536.585 ;
    RECT 0 536.655 0.070 536.725 ;
    RECT 0 536.795 0.070 536.865 ;
    RECT 0 536.935 0.070 537.005 ;
    RECT 0 537.075 0.070 537.145 ;
    RECT 0 537.215 0.070 537.285 ;
    RECT 0 537.355 0.070 537.425 ;
    RECT 0 537.495 0.070 537.565 ;
    RECT 0 537.635 0.070 537.705 ;
    RECT 0 537.775 0.070 537.845 ;
    RECT 0 537.915 0.070 537.985 ;
    RECT 0 538.055 0.070 538.125 ;
    RECT 0 538.195 0.070 538.265 ;
    RECT 0 538.335 0.070 538.405 ;
    RECT 0 538.475 0.070 538.545 ;
    RECT 0 538.615 0.070 538.685 ;
    RECT 0 538.755 0.070 538.825 ;
    RECT 0 538.895 0.070 538.965 ;
    RECT 0 539.035 0.070 539.105 ;
    RECT 0 539.175 0.070 539.245 ;
    RECT 0 539.315 0.070 539.385 ;
    RECT 0 539.455 0.070 539.525 ;
    RECT 0 539.595 0.070 539.665 ;
    RECT 0 539.735 0.070 539.805 ;
    RECT 0 539.875 0.070 539.945 ;
    RECT 0 540.015 0.070 540.085 ;
    RECT 0 540.155 0.070 540.225 ;
    RECT 0 540.295 0.070 540.365 ;
    RECT 0 540.435 0.070 540.505 ;
    RECT 0 540.575 0.070 540.645 ;
    RECT 0 540.715 0.070 540.785 ;
    RECT 0 540.855 0.070 540.925 ;
    RECT 0 540.995 0.070 541.065 ;
    RECT 0 541.135 0.070 541.205 ;
    RECT 0 541.275 0.070 541.345 ;
    RECT 0 541.415 0.070 541.485 ;
    RECT 0 541.555 0.070 541.625 ;
    RECT 0 541.695 0.070 541.765 ;
    RECT 0 541.835 0.070 541.905 ;
    RECT 0 541.975 0.070 542.045 ;
    RECT 0 542.115 0.070 542.185 ;
    RECT 0 542.255 0.070 542.325 ;
    RECT 0 542.395 0.070 542.465 ;
    RECT 0 542.535 0.070 542.605 ;
    RECT 0 542.675 0.070 542.745 ;
    RECT 0 542.815 0.070 542.885 ;
    RECT 0 542.955 0.070 543.025 ;
    RECT 0 543.095 0.070 543.165 ;
    RECT 0 543.235 0.070 543.305 ;
    RECT 0 543.375 0.070 543.445 ;
    RECT 0 543.515 0.070 543.585 ;
    RECT 0 543.655 0.070 543.725 ;
    RECT 0 543.795 0.070 543.865 ;
    RECT 0 543.935 0.070 544.005 ;
    RECT 0 544.075 0.070 544.145 ;
    RECT 0 544.215 0.070 544.285 ;
    RECT 0 544.355 0.070 544.425 ;
    RECT 0 544.495 0.070 544.565 ;
    RECT 0 544.635 0.070 544.705 ;
    RECT 0 544.775 0.070 544.845 ;
    RECT 0 544.915 0.070 544.985 ;
    RECT 0 545.055 0.070 545.125 ;
    RECT 0 545.195 0.070 545.265 ;
    RECT 0 545.335 0.070 545.405 ;
    RECT 0 545.475 0.070 545.545 ;
    RECT 0 545.615 0.070 545.685 ;
    RECT 0 545.755 0.070 545.825 ;
    RECT 0 545.895 0.070 545.965 ;
    RECT 0 546.035 0.070 546.105 ;
    RECT 0 546.175 0.070 546.245 ;
    RECT 0 546.315 0.070 546.385 ;
    RECT 0 546.455 0.070 546.525 ;
    RECT 0 546.595 0.070 546.665 ;
    RECT 0 546.735 0.070 546.805 ;
    RECT 0 546.875 0.070 546.945 ;
    RECT 0 547.015 0.070 547.085 ;
    RECT 0 547.155 0.070 547.225 ;
    RECT 0 547.295 0.070 547.365 ;
    RECT 0 547.435 0.070 547.505 ;
    RECT 0 547.575 0.070 547.645 ;
    RECT 0 547.715 0.070 547.785 ;
    RECT 0 547.855 0.070 547.925 ;
    RECT 0 547.995 0.070 548.065 ;
    RECT 0 548.135 0.070 548.205 ;
    RECT 0 548.275 0.070 548.345 ;
    RECT 0 548.415 0.070 548.485 ;
    RECT 0 548.555 0.070 548.625 ;
    RECT 0 548.695 0.070 548.765 ;
    RECT 0 548.835 0.070 548.905 ;
    RECT 0 548.975 0.070 549.045 ;
    RECT 0 549.115 0.070 549.185 ;
    RECT 0 549.255 0.070 549.325 ;
    RECT 0 549.395 0.070 549.465 ;
    RECT 0 549.535 0.070 549.605 ;
    RECT 0 549.675 0.070 549.745 ;
    RECT 0 549.815 0.070 549.885 ;
    RECT 0 549.955 0.070 550.025 ;
    RECT 0 550.095 0.070 550.165 ;
    RECT 0 550.235 0.070 550.305 ;
    RECT 0 550.375 0.070 550.445 ;
    RECT 0 550.515 0.070 550.585 ;
    RECT 0 550.655 0.070 550.725 ;
    RECT 0 550.795 0.070 550.865 ;
    RECT 0 550.935 0.070 551.005 ;
    RECT 0 551.075 0.070 551.145 ;
    RECT 0 551.215 0.070 551.285 ;
    RECT 0 551.355 0.070 551.425 ;
    RECT 0 551.495 0.070 551.565 ;
    RECT 0 551.635 0.070 551.705 ;
    RECT 0 551.775 0.070 551.845 ;
    RECT 0 551.915 0.070 551.985 ;
    RECT 0 552.055 0.070 552.125 ;
    RECT 0 552.195 0.070 552.265 ;
    RECT 0 552.335 0.070 552.405 ;
    RECT 0 552.475 0.070 552.545 ;
    RECT 0 552.615 0.070 552.685 ;
    RECT 0 552.755 0.070 552.825 ;
    RECT 0 552.895 0.070 552.965 ;
    RECT 0 553.035 0.070 553.105 ;
    RECT 0 553.175 0.070 553.245 ;
    RECT 0 553.315 0.070 553.385 ;
    RECT 0 553.455 0.070 553.525 ;
    RECT 0 553.595 0.070 553.665 ;
    RECT 0 553.735 0.070 553.805 ;
    RECT 0 553.875 0.070 553.945 ;
    RECT 0 554.015 0.070 554.085 ;
    RECT 0 554.155 0.070 554.225 ;
    RECT 0 554.295 0.070 554.365 ;
    RECT 0 554.435 0.070 554.505 ;
    RECT 0 554.575 0.070 554.645 ;
    RECT 0 554.715 0.070 554.785 ;
    RECT 0 554.855 0.070 554.925 ;
    RECT 0 554.995 0.070 555.065 ;
    RECT 0 555.135 0.070 555.205 ;
    RECT 0 555.275 0.070 555.345 ;
    RECT 0 555.415 0.070 555.485 ;
    RECT 0 555.555 0.070 555.625 ;
    RECT 0 555.695 0.070 555.765 ;
    RECT 0 555.835 0.070 555.905 ;
    RECT 0 555.975 0.070 556.045 ;
    RECT 0 556.115 0.070 556.185 ;
    RECT 0 556.255 0.070 556.325 ;
    RECT 0 556.395 0.070 556.465 ;
    RECT 0 556.535 0.070 556.605 ;
    RECT 0 556.675 0.070 556.745 ;
    RECT 0 556.815 0.070 556.885 ;
    RECT 0 556.955 0.070 557.025 ;
    RECT 0 557.095 0.070 557.165 ;
    RECT 0 557.235 0.070 557.305 ;
    RECT 0 557.375 0.070 557.445 ;
    RECT 0 557.515 0.070 557.585 ;
    RECT 0 557.655 0.070 557.725 ;
    RECT 0 557.795 0.070 557.865 ;
    RECT 0 557.935 0.070 558.005 ;
    RECT 0 558.075 0.070 558.145 ;
    RECT 0 558.215 0.070 558.285 ;
    RECT 0 558.355 0.070 558.425 ;
    RECT 0 558.495 0.070 558.565 ;
    RECT 0 558.635 0.070 558.705 ;
    RECT 0 558.775 0.070 558.845 ;
    RECT 0 558.915 0.070 558.985 ;
    RECT 0 559.055 0.070 559.125 ;
    RECT 0 559.195 0.070 559.265 ;
    RECT 0 559.335 0.070 559.405 ;
    RECT 0 559.475 0.070 559.545 ;
    RECT 0 559.615 0.070 559.685 ;
    RECT 0 559.755 0.070 559.825 ;
    RECT 0 559.895 0.070 559.965 ;
    RECT 0 560.035 0.070 560.105 ;
    RECT 0 560.175 0.070 560.245 ;
    RECT 0 560.315 0.070 560.385 ;
    RECT 0 560.455 0.070 560.525 ;
    RECT 0 560.595 0.070 560.665 ;
    RECT 0 560.735 0.070 560.805 ;
    RECT 0 560.875 0.070 560.945 ;
    RECT 0 561.015 0.070 561.085 ;
    RECT 0 561.155 0.070 561.225 ;
    RECT 0 561.295 0.070 561.365 ;
    RECT 0 561.435 0.070 561.505 ;
    RECT 0 561.575 0.070 561.645 ;
    RECT 0 561.715 0.070 561.785 ;
    RECT 0 561.855 0.070 561.925 ;
    RECT 0 561.995 0.070 562.065 ;
    RECT 0 562.135 0.070 562.205 ;
    RECT 0 562.275 0.070 562.345 ;
    RECT 0 562.415 0.070 562.485 ;
    RECT 0 562.555 0.070 562.625 ;
    RECT 0 562.695 0.070 562.765 ;
    RECT 0 562.835 0.070 562.905 ;
    RECT 0 562.975 0.070 563.045 ;
    RECT 0 563.115 0.070 563.185 ;
    RECT 0 563.255 0.070 563.325 ;
    RECT 0 563.395 0.070 563.465 ;
    RECT 0 563.535 0.070 563.605 ;
    RECT 0 563.675 0.070 563.745 ;
    RECT 0 563.815 0.070 563.885 ;
    RECT 0 563.955 0.070 564.025 ;
    RECT 0 564.095 0.070 564.165 ;
    RECT 0 564.235 0.070 564.305 ;
    RECT 0 564.375 0.070 564.445 ;
    RECT 0 564.515 0.070 564.585 ;
    RECT 0 564.655 0.070 564.725 ;
    RECT 0 564.795 0.070 564.865 ;
    RECT 0 564.935 0.070 565.005 ;
    RECT 0 565.075 0.070 565.145 ;
    RECT 0 565.215 0.070 565.285 ;
    RECT 0 565.355 0.070 565.425 ;
    RECT 0 565.495 0.070 565.565 ;
    RECT 0 565.635 0.070 565.705 ;
    RECT 0 565.775 0.070 565.845 ;
    RECT 0 565.915 0.070 565.985 ;
    RECT 0 566.055 0.070 566.125 ;
    RECT 0 566.195 0.070 566.265 ;
    RECT 0 566.335 0.070 566.405 ;
    RECT 0 566.475 0.070 566.545 ;
    RECT 0 566.615 0.070 566.685 ;
    RECT 0 566.755 0.070 566.825 ;
    RECT 0 566.895 0.070 566.965 ;
    RECT 0 567.035 0.070 567.105 ;
    RECT 0 567.175 0.070 567.245 ;
    RECT 0 567.315 0.070 567.385 ;
    RECT 0 567.455 0.070 567.525 ;
    RECT 0 567.595 0.070 567.665 ;
    RECT 0 567.735 0.070 567.805 ;
    RECT 0 567.875 0.070 567.945 ;
    RECT 0 568.015 0.070 568.085 ;
    RECT 0 568.155 0.070 568.225 ;
    RECT 0 568.295 0.070 568.365 ;
    RECT 0 568.435 0.070 568.505 ;
    RECT 0 568.575 0.070 568.645 ;
    RECT 0 568.715 0.070 568.785 ;
    RECT 0 568.855 0.070 568.925 ;
    RECT 0 568.995 0.070 569.065 ;
    RECT 0 569.135 0.070 569.205 ;
    RECT 0 569.275 0.070 569.345 ;
    RECT 0 569.415 0.070 569.485 ;
    RECT 0 569.555 0.070 569.625 ;
    RECT 0 569.695 0.070 569.765 ;
    RECT 0 569.835 0.070 569.905 ;
    RECT 0 569.975 0.070 570.045 ;
    RECT 0 570.115 0.070 570.185 ;
    RECT 0 570.255 0.070 570.325 ;
    RECT 0 570.395 0.070 570.465 ;
    RECT 0 570.535 0.070 570.605 ;
    RECT 0 570.675 0.070 570.745 ;
    RECT 0 570.815 0.070 570.885 ;
    RECT 0 570.955 0.070 571.025 ;
    RECT 0 571.095 0.070 571.165 ;
    RECT 0 571.235 0.070 571.305 ;
    RECT 0 571.375 0.070 571.445 ;
    RECT 0 571.515 0.070 571.585 ;
    RECT 0 571.655 0.070 571.725 ;
    RECT 0 571.795 0.070 571.865 ;
    RECT 0 571.935 0.070 572.005 ;
    RECT 0 572.075 0.070 572.145 ;
    RECT 0 572.215 0.070 572.285 ;
    RECT 0 572.355 0.070 572.425 ;
    RECT 0 572.495 0.070 572.565 ;
    RECT 0 572.635 0.070 572.705 ;
    RECT 0 572.775 0.070 572.845 ;
    RECT 0 572.915 0.070 572.985 ;
    RECT 0 573.055 0.070 573.125 ;
    RECT 0 573.195 0.070 573.265 ;
    RECT 0 573.335 0.070 573.405 ;
    RECT 0 573.475 0.070 573.545 ;
    RECT 0 573.615 0.070 573.685 ;
    RECT 0 573.755 0.070 573.825 ;
    RECT 0 573.895 0.070 573.965 ;
    RECT 0 574.035 0.070 574.105 ;
    RECT 0 574.175 0.070 574.245 ;
    RECT 0 574.315 0.070 574.385 ;
    RECT 0 574.455 0.070 574.525 ;
    RECT 0 574.595 0.070 574.665 ;
    RECT 0 574.735 0.070 574.805 ;
    RECT 0 574.875 0.070 574.945 ;
    RECT 0 575.015 0.070 575.085 ;
    RECT 0 575.155 0.070 575.225 ;
    RECT 0 575.295 0.070 575.365 ;
    RECT 0 575.435 0.070 575.505 ;
    RECT 0 575.575 0.070 575.645 ;
    RECT 0 575.715 0.070 575.785 ;
    RECT 0 575.855 0.070 575.925 ;
    RECT 0 575.995 0.070 576.065 ;
    RECT 0 576.135 0.070 576.205 ;
    RECT 0 576.275 0.070 576.345 ;
    RECT 0 576.415 0.070 576.485 ;
    RECT 0 576.555 0.070 576.625 ;
    RECT 0 576.695 0.070 576.765 ;
    RECT 0 576.835 0.070 576.905 ;
    RECT 0 576.975 0.070 577.045 ;
    RECT 0 577.115 0.070 577.185 ;
    RECT 0 577.255 0.070 577.325 ;
    RECT 0 577.395 0.070 577.465 ;
    RECT 0 577.535 0.070 577.605 ;
    RECT 0 577.675 0.070 577.745 ;
    RECT 0 577.815 0.070 577.885 ;
    RECT 0 577.955 0.070 578.025 ;
    RECT 0 578.095 0.070 578.165 ;
    RECT 0 578.235 0.070 578.305 ;
    RECT 0 578.375 0.070 578.445 ;
    RECT 0 578.515 0.070 578.585 ;
    RECT 0 578.655 0.070 578.725 ;
    RECT 0 578.795 0.070 578.865 ;
    RECT 0 578.935 0.070 579.005 ;
    RECT 0 579.075 0.070 579.145 ;
    RECT 0 579.215 0.070 579.285 ;
    RECT 0 579.355 0.070 579.425 ;
    RECT 0 579.495 0.070 579.565 ;
    RECT 0 579.635 0.070 579.705 ;
    RECT 0 579.775 0.070 579.845 ;
    RECT 0 579.915 0.070 579.985 ;
    RECT 0 580.055 0.070 580.125 ;
    RECT 0 580.195 0.070 580.265 ;
    RECT 0 580.335 0.070 580.405 ;
    RECT 0 580.475 0.070 580.545 ;
    RECT 0 580.615 0.070 580.685 ;
    RECT 0 580.755 0.070 580.825 ;
    RECT 0 580.895 0.070 580.965 ;
    RECT 0 581.035 0.070 581.105 ;
    RECT 0 581.175 0.070 581.245 ;
    RECT 0 581.315 0.070 581.385 ;
    RECT 0 581.455 0.070 581.525 ;
    RECT 0 581.595 0.070 581.665 ;
    RECT 0 581.735 0.070 581.805 ;
    RECT 0 581.875 0.070 581.945 ;
    RECT 0 582.015 0.070 582.085 ;
    RECT 0 582.155 0.070 582.225 ;
    RECT 0 582.295 0.070 582.365 ;
    RECT 0 582.435 0.070 582.505 ;
    RECT 0 582.575 0.070 582.645 ;
    RECT 0 582.715 0.070 582.785 ;
    RECT 0 582.855 0.070 582.925 ;
    RECT 0 582.995 0.070 583.065 ;
    RECT 0 583.135 0.070 583.205 ;
    RECT 0 583.275 0.070 583.345 ;
    RECT 0 583.415 0.070 583.485 ;
    RECT 0 583.555 0.070 583.625 ;
    RECT 0 583.695 0.070 583.765 ;
    RECT 0 583.835 0.070 583.905 ;
    RECT 0 583.975 0.070 584.045 ;
    RECT 0 584.115 0.070 584.185 ;
    RECT 0 584.255 0.070 584.325 ;
    RECT 0 584.395 0.070 584.465 ;
    RECT 0 584.535 0.070 584.605 ;
    RECT 0 584.675 0.070 584.745 ;
    RECT 0 584.815 0.070 584.885 ;
    RECT 0 584.955 0.070 585.025 ;
    RECT 0 585.095 0.070 585.165 ;
    RECT 0 585.235 0.070 585.305 ;
    RECT 0 585.375 0.070 585.445 ;
    RECT 0 585.515 0.070 585.585 ;
    RECT 0 585.655 0.070 585.725 ;
    RECT 0 585.795 0.070 585.865 ;
    RECT 0 585.935 0.070 586.005 ;
    RECT 0 586.075 0.070 586.145 ;
    RECT 0 586.215 0.070 586.285 ;
    RECT 0 586.355 0.070 586.425 ;
    RECT 0 586.495 0.070 586.565 ;
    RECT 0 586.635 0.070 586.705 ;
    RECT 0 586.775 0.070 586.845 ;
    RECT 0 586.915 0.070 586.985 ;
    RECT 0 587.055 0.070 587.125 ;
    RECT 0 587.195 0.070 587.265 ;
    RECT 0 587.335 0.070 587.405 ;
    RECT 0 587.475 0.070 587.545 ;
    RECT 0 587.615 0.070 587.685 ;
    RECT 0 587.755 0.070 587.825 ;
    RECT 0 587.895 0.070 587.965 ;
    RECT 0 588.035 0.070 588.105 ;
    RECT 0 588.175 0.070 588.245 ;
    RECT 0 588.315 0.070 588.385 ;
    RECT 0 588.455 0.070 588.525 ;
    RECT 0 588.595 0.070 588.665 ;
    RECT 0 588.735 0.070 588.805 ;
    RECT 0 588.875 0.070 588.945 ;
    RECT 0 589.015 0.070 589.085 ;
    RECT 0 589.155 0.070 589.225 ;
    RECT 0 589.295 0.070 589.365 ;
    RECT 0 589.435 0.070 589.505 ;
    RECT 0 589.575 0.070 589.645 ;
    RECT 0 589.715 0.070 589.785 ;
    RECT 0 589.855 0.070 589.925 ;
    RECT 0 589.995 0.070 590.065 ;
    RECT 0 590.135 0.070 590.205 ;
    RECT 0 590.275 0.070 590.345 ;
    RECT 0 590.415 0.070 590.485 ;
    RECT 0 590.555 0.070 590.625 ;
    RECT 0 590.695 0.070 590.765 ;
    RECT 0 590.835 0.070 590.905 ;
    RECT 0 590.975 0.070 591.045 ;
    RECT 0 591.115 0.070 591.185 ;
    RECT 0 591.255 0.070 591.325 ;
    RECT 0 591.395 0.070 591.465 ;
    RECT 0 591.535 0.070 591.605 ;
    RECT 0 591.675 0.070 591.745 ;
    RECT 0 591.815 0.070 591.885 ;
    RECT 0 591.955 0.070 592.025 ;
    RECT 0 592.095 0.070 592.165 ;
    RECT 0 592.235 0.070 592.305 ;
    RECT 0 592.375 0.070 592.445 ;
    RECT 0 592.515 0.070 592.585 ;
    RECT 0 592.655 0.070 592.725 ;
    RECT 0 592.795 0.070 592.865 ;
    RECT 0 592.935 0.070 593.005 ;
    RECT 0 593.075 0.070 593.145 ;
    RECT 0 593.215 0.070 593.285 ;
    RECT 0 593.355 0.070 593.425 ;
    RECT 0 593.495 0.070 593.565 ;
    RECT 0 593.635 0.070 593.705 ;
    RECT 0 593.775 0.070 593.845 ;
    RECT 0 593.915 0.070 593.985 ;
    RECT 0 594.055 0.070 594.125 ;
    RECT 0 594.195 0.070 594.265 ;
    RECT 0 594.335 0.070 594.405 ;
    RECT 0 594.475 0.070 594.545 ;
    RECT 0 594.615 0.070 594.685 ;
    RECT 0 594.755 0.070 594.825 ;
    RECT 0 594.895 0.070 594.965 ;
    RECT 0 595.035 0.070 595.105 ;
    RECT 0 595.175 0.070 595.245 ;
    RECT 0 595.315 0.070 595.385 ;
    RECT 0 595.455 0.070 595.525 ;
    RECT 0 595.595 0.070 595.665 ;
    RECT 0 595.735 0.070 595.805 ;
    RECT 0 595.875 0.070 595.945 ;
    RECT 0 596.015 0.070 596.085 ;
    RECT 0 596.155 0.070 596.225 ;
    RECT 0 596.295 0.070 596.365 ;
    RECT 0 596.435 0.070 596.505 ;
    RECT 0 596.575 0.070 596.645 ;
    RECT 0 596.715 0.070 596.785 ;
    RECT 0 596.855 0.070 596.925 ;
    RECT 0 596.995 0.070 597.065 ;
    RECT 0 597.135 0.070 597.205 ;
    RECT 0 597.275 0.070 597.345 ;
    RECT 0 597.415 0.070 597.485 ;
    RECT 0 597.555 0.070 597.625 ;
    RECT 0 597.695 0.070 597.765 ;
    RECT 0 597.835 0.070 597.905 ;
    RECT 0 597.975 0.070 598.045 ;
    RECT 0 598.115 0.070 598.185 ;
    RECT 0 598.255 0.070 598.325 ;
    RECT 0 598.395 0.070 598.465 ;
    RECT 0 598.535 0.070 598.605 ;
    RECT 0 598.675 0.070 598.745 ;
    RECT 0 598.815 0.070 598.885 ;
    RECT 0 598.955 0.070 599.025 ;
    RECT 0 599.095 0.070 599.165 ;
    RECT 0 599.235 0.070 599.305 ;
    RECT 0 599.375 0.070 599.445 ;
    RECT 0 599.515 0.070 599.585 ;
    RECT 0 599.655 0.070 599.725 ;
    RECT 0 599.795 0.070 599.865 ;
    RECT 0 599.935 0.070 600.005 ;
    RECT 0 600.075 0.070 600.145 ;
    RECT 0 600.215 0.070 600.285 ;
    RECT 0 600.355 0.070 600.425 ;
    RECT 0 600.495 0.070 600.565 ;
    RECT 0 600.635 0.070 600.705 ;
    RECT 0 600.775 0.070 600.845 ;
    RECT 0 600.915 0.070 600.985 ;
    RECT 0 601.055 0.070 601.125 ;
    RECT 0 601.195 0.070 601.265 ;
    RECT 0 601.335 0.070 601.405 ;
    RECT 0 601.475 0.070 601.545 ;
    RECT 0 601.615 0.070 601.685 ;
    RECT 0 601.755 0.070 601.825 ;
    RECT 0 601.895 0.070 601.965 ;
    RECT 0 602.035 0.070 602.105 ;
    RECT 0 602.175 0.070 602.245 ;
    RECT 0 602.315 0.070 602.385 ;
    RECT 0 602.455 0.070 602.525 ;
    RECT 0 602.595 0.070 602.665 ;
    RECT 0 602.735 0.070 602.805 ;
    RECT 0 602.875 0.070 602.945 ;
    RECT 0 603.015 0.070 603.085 ;
    RECT 0 603.155 0.070 603.225 ;
    RECT 0 603.295 0.070 603.365 ;
    RECT 0 603.435 0.070 603.505 ;
    RECT 0 603.575 0.070 603.645 ;
    RECT 0 603.715 0.070 603.785 ;
    RECT 0 603.855 0.070 603.925 ;
    RECT 0 603.995 0.070 604.065 ;
    RECT 0 604.135 0.070 604.205 ;
    RECT 0 604.275 0.070 604.345 ;
    RECT 0 604.415 0.070 604.485 ;
    RECT 0 604.555 0.070 604.625 ;
    RECT 0 604.695 0.070 604.765 ;
    RECT 0 604.835 0.070 604.905 ;
    RECT 0 604.975 0.070 605.045 ;
    RECT 0 605.115 0.070 605.185 ;
    RECT 0 605.255 0.070 605.325 ;
    RECT 0 605.395 0.070 605.465 ;
    RECT 0 605.535 0.070 605.605 ;
    RECT 0 605.675 0.070 605.745 ;
    RECT 0 605.815 0.070 605.885 ;
    RECT 0 605.955 0.070 606.025 ;
    RECT 0 606.095 0.070 606.165 ;
    RECT 0 606.235 0.070 606.305 ;
    RECT 0 606.375 0.070 606.445 ;
    RECT 0 606.515 0.070 606.585 ;
    RECT 0 606.655 0.070 606.725 ;
    RECT 0 606.795 0.070 606.865 ;
    RECT 0 606.935 0.070 607.005 ;
    RECT 0 607.075 0.070 607.145 ;
    RECT 0 607.215 0.070 607.285 ;
    RECT 0 607.355 0.070 607.425 ;
    RECT 0 607.495 0.070 607.565 ;
    RECT 0 607.635 0.070 607.705 ;
    RECT 0 607.775 0.070 607.845 ;
    RECT 0 607.915 0.070 607.985 ;
    RECT 0 608.055 0.070 608.125 ;
    RECT 0 608.195 0.070 608.265 ;
    RECT 0 608.335 0.070 608.405 ;
    RECT 0 608.475 0.070 608.545 ;
    RECT 0 608.615 0.070 608.685 ;
    RECT 0 608.755 0.070 608.825 ;
    RECT 0 608.895 0.070 608.965 ;
    RECT 0 609.035 0.070 609.105 ;
    RECT 0 609.175 0.070 609.245 ;
    RECT 0 609.315 0.070 609.385 ;
    RECT 0 609.455 0.070 609.525 ;
    RECT 0 609.595 0.070 609.665 ;
    RECT 0 609.735 0.070 609.805 ;
    RECT 0 609.875 0.070 609.945 ;
    RECT 0 610.015 0.070 610.085 ;
    RECT 0 610.155 0.070 610.225 ;
    RECT 0 610.295 0.070 610.365 ;
    RECT 0 610.435 0.070 610.505 ;
    RECT 0 610.575 0.070 610.645 ;
    RECT 0 610.715 0.070 610.785 ;
    RECT 0 610.855 0.070 610.925 ;
    RECT 0 610.995 0.070 611.065 ;
    RECT 0 611.135 0.070 611.205 ;
    RECT 0 611.275 0.070 611.345 ;
    RECT 0 611.415 0.070 611.485 ;
    RECT 0 611.555 0.070 611.625 ;
    RECT 0 611.695 0.070 611.765 ;
    RECT 0 611.835 0.070 611.905 ;
    RECT 0 611.975 0.070 612.045 ;
    RECT 0 612.115 0.070 612.185 ;
    RECT 0 612.255 0.070 612.325 ;
    RECT 0 612.395 0.070 612.465 ;
    RECT 0 612.535 0.070 612.605 ;
    RECT 0 612.675 0.070 612.745 ;
    RECT 0 612.815 0.070 612.885 ;
    RECT 0 612.955 0.070 613.025 ;
    RECT 0 613.095 0.070 613.165 ;
    RECT 0 613.235 0.070 613.305 ;
    RECT 0 613.375 0.070 613.445 ;
    RECT 0 613.515 0.070 613.585 ;
    RECT 0 613.655 0.070 613.725 ;
    RECT 0 613.795 0.070 613.865 ;
    RECT 0 613.935 0.070 614.005 ;
    RECT 0 614.075 0.070 614.145 ;
    RECT 0 614.215 0.070 614.285 ;
    RECT 0 614.355 0.070 614.425 ;
    RECT 0 614.495 0.070 614.565 ;
    RECT 0 614.635 0.070 614.705 ;
    RECT 0 614.775 0.070 614.845 ;
    RECT 0 614.915 0.070 614.985 ;
    RECT 0 615.055 0.070 615.125 ;
    RECT 0 615.195 0.070 615.265 ;
    RECT 0 615.335 0.070 615.405 ;
    RECT 0 615.475 0.070 615.545 ;
    RECT 0 615.615 0.070 615.685 ;
    RECT 0 615.755 0.070 615.825 ;
    RECT 0 615.895 0.070 615.965 ;
    RECT 0 616.035 0.070 616.105 ;
    RECT 0 616.175 0.070 616.245 ;
    RECT 0 616.315 0.070 616.385 ;
    RECT 0 616.455 0.070 616.525 ;
    RECT 0 616.595 0.070 616.665 ;
    RECT 0 616.735 0.070 616.805 ;
    RECT 0 616.875 0.070 616.945 ;
    RECT 0 617.015 0.070 617.085 ;
    RECT 0 617.155 0.070 617.225 ;
    RECT 0 617.295 0.070 617.365 ;
    RECT 0 617.435 0.070 617.505 ;
    RECT 0 617.575 0.070 617.645 ;
    RECT 0 617.715 0.070 617.785 ;
    RECT 0 617.855 0.070 617.925 ;
    RECT 0 617.995 0.070 618.065 ;
    RECT 0 618.135 0.070 618.205 ;
    RECT 0 618.275 0.070 618.345 ;
    RECT 0 618.415 0.070 618.485 ;
    RECT 0 618.555 0.070 618.625 ;
    RECT 0 618.695 0.070 618.765 ;
    RECT 0 618.835 0.070 618.905 ;
    RECT 0 618.975 0.070 619.045 ;
    RECT 0 619.115 0.070 619.185 ;
    RECT 0 619.255 0.070 619.325 ;
    RECT 0 619.395 0.070 619.465 ;
    RECT 0 619.535 0.070 619.605 ;
    RECT 0 619.675 0.070 619.745 ;
    RECT 0 619.815 0.070 619.885 ;
    RECT 0 619.955 0.070 620.025 ;
    RECT 0 620.095 0.070 620.165 ;
    RECT 0 620.235 0.070 620.305 ;
    RECT 0 620.375 0.070 620.445 ;
    RECT 0 620.515 0.070 620.585 ;
    RECT 0 620.655 0.070 620.725 ;
    RECT 0 620.795 0.070 620.865 ;
    RECT 0 620.935 0.070 621.005 ;
    RECT 0 621.075 0.070 621.145 ;
    RECT 0 621.215 0.070 621.285 ;
    RECT 0 621.355 0.070 621.425 ;
    RECT 0 621.495 0.070 621.565 ;
    RECT 0 621.635 0.070 621.705 ;
    RECT 0 621.775 0.070 621.845 ;
    RECT 0 621.915 0.070 621.985 ;
    RECT 0 622.055 0.070 622.125 ;
    RECT 0 622.195 0.070 622.265 ;
    RECT 0 622.335 0.070 622.405 ;
    RECT 0 622.475 0.070 622.545 ;
    RECT 0 622.615 0.070 622.685 ;
    RECT 0 622.755 0.070 622.825 ;
    RECT 0 622.895 0.070 622.965 ;
    RECT 0 623.035 0.070 623.105 ;
    RECT 0 623.175 0.070 623.245 ;
    RECT 0 623.315 0.070 623.385 ;
    RECT 0 623.455 0.070 623.525 ;
    RECT 0 623.595 0.070 623.665 ;
    RECT 0 623.735 0.070 623.805 ;
    RECT 0 623.875 0.070 623.945 ;
    RECT 0 624.015 0.070 624.085 ;
    RECT 0 624.155 0.070 624.225 ;
    RECT 0 624.295 0.070 624.365 ;
    RECT 0 624.435 0.070 624.505 ;
    RECT 0 624.575 0.070 624.645 ;
    RECT 0 624.715 0.070 624.785 ;
    RECT 0 624.855 0.070 624.925 ;
    RECT 0 624.995 0.070 625.065 ;
    RECT 0 625.135 0.070 625.205 ;
    RECT 0 625.275 0.070 625.345 ;
    RECT 0 625.415 0.070 625.485 ;
    RECT 0 625.555 0.070 625.625 ;
    RECT 0 625.695 0.070 625.765 ;
    RECT 0 625.835 0.070 625.905 ;
    RECT 0 625.975 0.070 626.045 ;
    RECT 0 626.115 0.070 626.185 ;
    RECT 0 626.255 0.070 626.325 ;
    RECT 0 626.395 0.070 626.465 ;
    RECT 0 626.535 0.070 626.605 ;
    RECT 0 626.675 0.070 626.745 ;
    RECT 0 626.815 0.070 626.885 ;
    RECT 0 626.955 0.070 627.025 ;
    RECT 0 627.095 0.070 627.165 ;
    RECT 0 627.235 0.070 627.305 ;
    RECT 0 627.375 0.070 627.445 ;
    RECT 0 627.515 0.070 627.585 ;
    RECT 0 627.655 0.070 627.725 ;
    RECT 0 627.795 0.070 627.865 ;
    RECT 0 627.935 0.070 628.005 ;
    RECT 0 628.075 0.070 628.145 ;
    RECT 0 628.215 0.070 628.285 ;
    RECT 0 628.355 0.070 628.425 ;
    RECT 0 628.495 0.070 628.565 ;
    RECT 0 628.635 0.070 628.705 ;
    RECT 0 628.775 0.070 628.845 ;
    RECT 0 628.915 0.070 628.985 ;
    RECT 0 629.055 0.070 629.125 ;
    RECT 0 629.195 0.070 629.265 ;
    RECT 0 629.335 0.070 629.405 ;
    RECT 0 629.475 0.070 629.545 ;
    RECT 0 629.615 0.070 629.685 ;
    RECT 0 629.755 0.070 629.825 ;
    RECT 0 629.895 0.070 629.965 ;
    RECT 0 630.035 0.070 630.105 ;
    RECT 0 630.175 0.070 630.245 ;
    RECT 0 630.315 0.070 630.385 ;
    RECT 0 630.455 0.070 630.525 ;
    RECT 0 630.595 0.070 630.665 ;
    RECT 0 630.735 0.070 630.805 ;
    RECT 0 630.875 0.070 630.945 ;
    RECT 0 631.015 0.070 631.085 ;
    RECT 0 631.155 0.070 631.225 ;
    RECT 0 631.295 0.070 631.365 ;
    RECT 0 631.435 0.070 631.505 ;
    RECT 0 631.575 0.070 631.645 ;
    RECT 0 631.715 0.070 631.785 ;
    RECT 0 631.855 0.070 631.925 ;
    RECT 0 631.995 0.070 632.065 ;
    RECT 0 632.135 0.070 632.205 ;
    RECT 0 632.275 0.070 632.345 ;
    RECT 0 632.415 0.070 632.485 ;
    RECT 0 632.555 0.070 632.625 ;
    RECT 0 632.695 0.070 632.765 ;
    RECT 0 632.835 0.070 632.905 ;
    RECT 0 632.975 0.070 633.045 ;
    RECT 0 633.115 0.070 633.185 ;
    RECT 0 633.255 0.070 633.325 ;
    RECT 0 633.395 0.070 633.465 ;
    RECT 0 633.535 0.070 633.605 ;
    RECT 0 633.675 0.070 633.745 ;
    RECT 0 633.815 0.070 633.885 ;
    RECT 0 633.955 0.070 634.025 ;
    RECT 0 634.095 0.070 634.165 ;
    RECT 0 634.235 0.070 634.305 ;
    RECT 0 634.375 0.070 634.445 ;
    RECT 0 634.515 0.070 634.585 ;
    RECT 0 634.655 0.070 634.725 ;
    RECT 0 634.795 0.070 634.865 ;
    RECT 0 634.935 0.070 635.005 ;
    RECT 0 635.075 0.070 635.145 ;
    RECT 0 635.215 0.070 635.285 ;
    RECT 0 635.355 0.070 635.425 ;
    RECT 0 635.495 0.070 635.565 ;
    RECT 0 635.635 0.070 635.705 ;
    RECT 0 635.775 0.070 635.845 ;
    RECT 0 635.915 0.070 635.985 ;
    RECT 0 636.055 0.070 636.125 ;
    RECT 0 636.195 0.070 636.265 ;
    RECT 0 636.335 0.070 636.405 ;
    RECT 0 636.475 0.070 636.545 ;
    RECT 0 636.615 0.070 636.685 ;
    RECT 0 636.755 0.070 636.825 ;
    RECT 0 636.895 0.070 636.965 ;
    RECT 0 637.035 0.070 637.105 ;
    RECT 0 637.175 0.070 637.245 ;
    RECT 0 637.315 0.070 637.385 ;
    RECT 0 637.455 0.070 637.525 ;
    RECT 0 637.595 0.070 637.665 ;
    RECT 0 637.735 0.070 637.805 ;
    RECT 0 637.875 0.070 637.945 ;
    RECT 0 638.015 0.070 638.085 ;
    RECT 0 638.155 0.070 638.225 ;
    RECT 0 638.295 0.070 638.365 ;
    RECT 0 638.435 0.070 638.505 ;
    RECT 0 638.575 0.070 638.645 ;
    RECT 0 638.715 0.070 638.785 ;
    RECT 0 638.855 0.070 638.925 ;
    RECT 0 638.995 0.070 639.065 ;
    RECT 0 639.135 0.070 639.205 ;
    RECT 0 639.275 0.070 639.345 ;
    RECT 0 639.415 0.070 639.485 ;
    RECT 0 639.555 0.070 639.625 ;
    RECT 0 639.695 0.070 639.765 ;
    RECT 0 639.835 0.070 639.905 ;
    RECT 0 639.975 0.070 640.045 ;
    RECT 0 640.115 0.070 640.185 ;
    RECT 0 640.255 0.070 640.325 ;
    RECT 0 640.395 0.070 640.465 ;
    RECT 0 640.535 0.070 640.605 ;
    RECT 0 640.675 0.070 640.745 ;
    RECT 0 640.815 0.070 640.885 ;
    RECT 0 640.955 0.070 641.025 ;
    RECT 0 641.095 0.070 641.165 ;
    RECT 0 641.235 0.070 641.305 ;
    RECT 0 641.375 0.070 641.445 ;
    RECT 0 641.515 0.070 641.585 ;
    RECT 0 641.655 0.070 641.725 ;
    RECT 0 641.795 0.070 641.865 ;
    RECT 0 641.935 0.070 642.005 ;
    RECT 0 642.075 0.070 642.145 ;
    RECT 0 642.215 0.070 642.285 ;
    RECT 0 642.355 0.070 642.425 ;
    RECT 0 642.495 0.070 642.565 ;
    RECT 0 642.635 0.070 642.705 ;
    RECT 0 642.775 0.070 642.845 ;
    RECT 0 642.915 0.070 642.985 ;
    RECT 0 643.055 0.070 643.125 ;
    RECT 0 643.195 0.070 643.265 ;
    RECT 0 643.335 0.070 643.405 ;
    RECT 0 643.475 0.070 643.545 ;
    RECT 0 643.615 0.070 643.685 ;
    RECT 0 643.755 0.070 643.825 ;
    RECT 0 643.895 0.070 643.965 ;
    RECT 0 644.035 0.070 644.105 ;
    RECT 0 644.175 0.070 644.245 ;
    RECT 0 644.315 0.070 644.385 ;
    RECT 0 644.455 0.070 644.525 ;
    RECT 0 644.595 0.070 644.665 ;
    RECT 0 644.735 0.070 644.805 ;
    RECT 0 644.875 0.070 644.945 ;
    RECT 0 645.015 0.070 645.085 ;
    RECT 0 645.155 0.070 645.225 ;
    RECT 0 645.295 0.070 645.365 ;
    RECT 0 645.435 0.070 645.505 ;
    RECT 0 645.575 0.070 645.645 ;
    RECT 0 645.715 0.070 645.785 ;
    RECT 0 645.855 0.070 645.925 ;
    RECT 0 645.995 0.070 646.065 ;
    RECT 0 646.135 0.070 646.205 ;
    RECT 0 646.275 0.070 646.345 ;
    RECT 0 646.415 0.070 646.485 ;
    RECT 0 646.555 0.070 646.625 ;
    RECT 0 646.695 0.070 646.765 ;
    RECT 0 646.835 0.070 646.905 ;
    RECT 0 646.975 0.070 647.045 ;
    RECT 0 647.115 0.070 647.185 ;
    RECT 0 647.255 0.070 647.325 ;
    RECT 0 647.395 0.070 647.465 ;
    RECT 0 647.535 0.070 647.605 ;
    RECT 0 647.675 0.070 647.745 ;
    RECT 0 647.815 0.070 647.885 ;
    RECT 0 647.955 0.070 648.025 ;
    RECT 0 648.095 0.070 648.165 ;
    RECT 0 648.235 0.070 648.305 ;
    RECT 0 648.375 0.070 648.445 ;
    RECT 0 648.515 0.070 648.585 ;
    RECT 0 648.655 0.070 648.725 ;
    RECT 0 648.795 0.070 648.865 ;
    RECT 0 648.935 0.070 649.005 ;
    RECT 0 649.075 0.070 649.145 ;
    RECT 0 649.215 0.070 649.285 ;
    RECT 0 649.355 0.070 649.425 ;
    RECT 0 649.495 0.070 649.565 ;
    RECT 0 649.635 0.070 649.705 ;
    RECT 0 649.775 0.070 649.845 ;
    RECT 0 649.915 0.070 649.985 ;
    RECT 0 650.055 0.070 650.125 ;
    RECT 0 650.195 0.070 650.265 ;
    RECT 0 650.335 0.070 650.405 ;
    RECT 0 650.475 0.070 650.545 ;
    RECT 0 650.615 0.070 650.685 ;
    RECT 0 650.755 0.070 650.825 ;
    RECT 0 650.895 0.070 650.965 ;
    RECT 0 651.035 0.070 651.105 ;
    RECT 0 651.175 0.070 651.245 ;
    RECT 0 651.315 0.070 651.385 ;
    RECT 0 651.455 0.070 651.525 ;
    RECT 0 651.595 0.070 651.665 ;
    RECT 0 651.735 0.070 651.805 ;
    RECT 0 651.875 0.070 651.945 ;
    RECT 0 652.015 0.070 652.085 ;
    RECT 0 652.155 0.070 652.225 ;
    RECT 0 652.295 0.070 652.365 ;
    RECT 0 652.435 0.070 652.505 ;
    RECT 0 652.575 0.070 652.645 ;
    RECT 0 652.715 0.070 652.785 ;
    RECT 0 652.855 0.070 652.925 ;
    RECT 0 652.995 0.070 653.065 ;
    RECT 0 653.135 0.070 653.205 ;
    RECT 0 653.275 0.070 653.345 ;
    RECT 0 653.415 0.070 653.485 ;
    RECT 0 653.555 0.070 653.625 ;
    RECT 0 653.695 0.070 653.765 ;
    RECT 0 653.835 0.070 653.905 ;
    RECT 0 653.975 0.070 654.045 ;
    RECT 0 654.115 0.070 654.185 ;
    RECT 0 654.255 0.070 654.325 ;
    RECT 0 654.395 0.070 654.465 ;
    RECT 0 654.535 0.070 654.605 ;
    RECT 0 654.675 0.070 654.745 ;
    RECT 0 654.815 0.070 654.885 ;
    RECT 0 654.955 0.070 655.025 ;
    RECT 0 655.095 0.070 655.165 ;
    RECT 0 655.235 0.070 655.305 ;
    RECT 0 655.375 0.070 655.445 ;
    RECT 0 655.515 0.070 655.585 ;
    RECT 0 655.655 0.070 655.725 ;
    RECT 0 655.795 0.070 655.865 ;
    RECT 0 655.935 0.070 656.005 ;
    RECT 0 656.075 0.070 656.145 ;
    RECT 0 656.215 0.070 656.285 ;
    RECT 0 656.355 0.070 656.425 ;
    RECT 0 656.495 0.070 656.565 ;
    RECT 0 656.635 0.070 656.705 ;
    RECT 0 656.775 0.070 656.845 ;
    RECT 0 656.915 0.070 656.985 ;
    RECT 0 657.055 0.070 657.125 ;
    RECT 0 657.195 0.070 657.265 ;
    RECT 0 657.335 0.070 657.405 ;
    RECT 0 657.475 0.070 657.545 ;
    RECT 0 657.615 0.070 657.685 ;
    RECT 0 657.755 0.070 657.825 ;
    RECT 0 657.895 0.070 657.965 ;
    RECT 0 658.035 0.070 658.105 ;
    RECT 0 658.175 0.070 658.245 ;
    RECT 0 658.315 0.070 658.385 ;
    RECT 0 658.455 0.070 658.525 ;
    RECT 0 658.595 0.070 658.665 ;
    RECT 0 658.735 0.070 658.805 ;
    RECT 0 658.875 0.070 658.945 ;
    RECT 0 659.015 0.070 659.085 ;
    RECT 0 659.155 0.070 659.225 ;
    RECT 0 659.295 0.070 659.365 ;
    RECT 0 659.435 0.070 659.505 ;
    RECT 0 659.575 0.070 659.645 ;
    RECT 0 659.715 0.070 659.785 ;
    RECT 0 659.855 0.070 659.925 ;
    RECT 0 659.995 0.070 660.065 ;
    RECT 0 660.135 0.070 660.205 ;
    RECT 0 660.275 0.070 660.345 ;
    RECT 0 660.415 0.070 660.485 ;
    RECT 0 660.555 0.070 660.625 ;
    RECT 0 660.695 0.070 660.765 ;
    RECT 0 660.835 0.070 660.905 ;
    RECT 0 660.975 0.070 661.045 ;
    RECT 0 661.115 0.070 661.185 ;
    RECT 0 661.255 0.070 661.325 ;
    RECT 0 661.395 0.070 661.465 ;
    RECT 0 661.535 0.070 661.605 ;
    RECT 0 661.675 0.070 661.745 ;
    RECT 0 661.815 0.070 661.885 ;
    RECT 0 661.955 0.070 662.025 ;
    RECT 0 662.095 0.070 662.165 ;
    RECT 0 662.235 0.070 662.305 ;
    RECT 0 662.375 0.070 662.445 ;
    RECT 0 662.515 0.070 662.585 ;
    RECT 0 662.655 0.070 662.725 ;
    RECT 0 662.795 0.070 662.865 ;
    RECT 0 662.935 0.070 663.005 ;
    RECT 0 663.075 0.070 663.145 ;
    RECT 0 663.215 0.070 663.285 ;
    RECT 0 663.355 0.070 663.425 ;
    RECT 0 663.495 0.070 663.565 ;
    RECT 0 663.635 0.070 663.705 ;
    RECT 0 663.775 0.070 663.845 ;
    RECT 0 663.915 0.070 663.985 ;
    RECT 0 664.055 0.070 664.125 ;
    RECT 0 664.195 0.070 664.265 ;
    RECT 0 664.335 0.070 664.405 ;
    RECT 0 664.475 0.070 664.545 ;
    RECT 0 664.615 0.070 664.685 ;
    RECT 0 664.755 0.070 664.825 ;
    RECT 0 664.895 0.070 664.965 ;
    RECT 0 665.035 0.070 665.105 ;
    RECT 0 665.175 0.070 665.245 ;
    RECT 0 665.315 0.070 665.385 ;
    RECT 0 665.455 0.070 665.525 ;
    RECT 0 665.595 0.070 665.665 ;
    RECT 0 665.735 0.070 665.805 ;
    RECT 0 665.875 0.070 665.945 ;
    RECT 0 666.015 0.070 666.085 ;
    RECT 0 666.155 0.070 666.225 ;
    RECT 0 666.295 0.070 666.365 ;
    RECT 0 666.435 0.070 666.505 ;
    RECT 0 666.575 0.070 666.645 ;
    RECT 0 666.715 0.070 666.785 ;
    RECT 0 666.855 0.070 666.925 ;
    RECT 0 666.995 0.070 667.065 ;
    RECT 0 667.135 0.070 667.205 ;
    RECT 0 667.275 0.070 667.345 ;
    RECT 0 667.415 0.070 667.485 ;
    RECT 0 667.555 0.070 667.625 ;
    RECT 0 667.695 0.070 667.765 ;
    RECT 0 667.835 0.070 667.905 ;
    RECT 0 667.975 0.070 668.045 ;
    RECT 0 668.115 0.070 668.185 ;
    RECT 0 668.255 0.070 668.325 ;
    RECT 0 668.395 0.070 668.465 ;
    RECT 0 668.535 0.070 668.605 ;
    RECT 0 668.675 0.070 668.745 ;
    RECT 0 668.815 0.070 668.885 ;
    RECT 0 668.955 0.070 669.025 ;
    RECT 0 669.095 0.070 669.165 ;
    RECT 0 669.235 0.070 669.305 ;
    RECT 0 669.375 0.070 669.445 ;
    RECT 0 669.515 0.070 669.585 ;
    RECT 0 669.655 0.070 669.725 ;
    RECT 0 669.795 0.070 669.865 ;
    RECT 0 669.935 0.070 670.005 ;
    RECT 0 670.075 0.070 670.145 ;
    RECT 0 670.215 0.070 670.285 ;
    RECT 0 670.355 0.070 670.425 ;
    RECT 0 670.495 0.070 670.565 ;
    RECT 0 670.635 0.070 670.705 ;
    RECT 0 670.775 0.070 670.845 ;
    RECT 0 670.915 0.070 670.985 ;
    RECT 0 671.055 0.070 671.125 ;
    RECT 0 671.195 0.070 671.265 ;
    RECT 0 671.335 0.070 671.405 ;
    RECT 0 671.475 0.070 671.545 ;
    RECT 0 671.615 0.070 671.685 ;
    RECT 0 671.755 0.070 671.825 ;
    RECT 0 671.895 0.070 671.965 ;
    RECT 0 672.035 0.070 672.105 ;
    RECT 0 672.175 0.070 672.245 ;
    RECT 0 672.315 0.070 672.385 ;
    RECT 0 672.455 0.070 672.525 ;
    RECT 0 672.595 0.070 672.665 ;
    RECT 0 672.735 0.070 672.805 ;
    RECT 0 672.875 0.070 672.945 ;
    RECT 0 673.015 0.070 673.085 ;
    RECT 0 673.155 0.070 673.225 ;
    RECT 0 673.295 0.070 673.365 ;
    RECT 0 673.435 0.070 673.505 ;
    RECT 0 673.575 0.070 673.645 ;
    RECT 0 673.715 0.070 673.785 ;
    RECT 0 673.855 0.070 673.925 ;
    RECT 0 673.995 0.070 674.065 ;
    RECT 0 674.135 0.070 674.205 ;
    RECT 0 674.275 0.070 674.345 ;
    RECT 0 674.415 0.070 674.485 ;
    RECT 0 674.555 0.070 674.625 ;
    RECT 0 674.695 0.070 674.765 ;
    RECT 0 674.835 0.070 674.905 ;
    RECT 0 674.975 0.070 675.045 ;
    RECT 0 675.115 0.070 675.185 ;
    RECT 0 675.255 0.070 675.325 ;
    RECT 0 675.395 0.070 675.465 ;
    RECT 0 675.535 0.070 675.605 ;
    RECT 0 675.675 0.070 675.745 ;
    RECT 0 675.815 0.070 675.885 ;
    RECT 0 675.955 0.070 676.025 ;
    RECT 0 676.095 0.070 676.165 ;
    RECT 0 676.235 0.070 676.305 ;
    RECT 0 676.375 0.070 676.445 ;
    RECT 0 676.515 0.070 676.585 ;
    RECT 0 676.655 0.070 676.725 ;
    RECT 0 676.795 0.070 676.865 ;
    RECT 0 676.935 0.070 677.005 ;
    RECT 0 677.075 0.070 677.145 ;
    RECT 0 677.215 0.070 677.285 ;
    RECT 0 677.355 0.070 677.425 ;
    RECT 0 677.495 0.070 677.565 ;
    RECT 0 677.635 0.070 677.705 ;
    RECT 0 677.775 0.070 677.845 ;
    RECT 0 677.915 0.070 677.985 ;
    RECT 0 678.055 0.070 678.125 ;
    RECT 0 678.195 0.070 678.265 ;
    RECT 0 678.335 0.070 678.405 ;
    RECT 0 678.475 0.070 678.545 ;
    RECT 0 678.615 0.070 678.685 ;
    RECT 0 678.755 0.070 678.825 ;
    RECT 0 678.895 0.070 678.965 ;
    RECT 0 679.035 0.070 679.105 ;
    RECT 0 679.175 0.070 679.245 ;
    RECT 0 679.315 0.070 679.385 ;
    RECT 0 679.455 0.070 679.525 ;
    RECT 0 679.595 0.070 679.665 ;
    RECT 0 679.735 0.070 679.805 ;
    RECT 0 679.875 0.070 679.945 ;
    RECT 0 680.015 0.070 680.085 ;
    RECT 0 680.155 0.070 680.225 ;
    RECT 0 680.295 0.070 680.365 ;
    RECT 0 680.435 0.070 680.505 ;
    RECT 0 680.575 0.070 680.645 ;
    RECT 0 680.715 0.070 680.785 ;
    RECT 0 680.855 0.070 680.925 ;
    RECT 0 680.995 0.070 681.065 ;
    RECT 0 681.135 0.070 681.205 ;
    RECT 0 681.275 0.070 681.345 ;
    RECT 0 681.415 0.070 681.485 ;
    RECT 0 681.555 0.070 681.625 ;
    RECT 0 681.695 0.070 681.765 ;
    RECT 0 681.835 0.070 681.905 ;
    RECT 0 681.975 0.070 682.045 ;
    RECT 0 682.115 0.070 682.185 ;
    RECT 0 682.255 0.070 682.325 ;
    RECT 0 682.395 0.070 682.465 ;
    RECT 0 682.535 0.070 682.605 ;
    RECT 0 682.675 0.070 682.745 ;
    RECT 0 682.815 0.070 682.885 ;
    RECT 0 682.955 0.070 683.025 ;
    RECT 0 683.095 0.070 683.165 ;
    RECT 0 683.235 0.070 683.305 ;
    RECT 0 683.375 0.070 683.445 ;
    RECT 0 683.515 0.070 683.585 ;
    RECT 0 683.655 0.070 683.725 ;
    RECT 0 683.795 0.070 683.865 ;
    RECT 0 683.935 0.070 684.005 ;
    RECT 0 684.075 0.070 684.145 ;
    RECT 0 684.215 0.070 684.285 ;
    RECT 0 684.355 0.070 684.425 ;
    RECT 0 684.495 0.070 684.565 ;
    RECT 0 684.635 0.070 684.705 ;
    RECT 0 684.775 0.070 684.845 ;
    RECT 0 684.915 0.070 684.985 ;
    RECT 0 685.055 0.070 685.125 ;
    RECT 0 685.195 0.070 685.265 ;
    RECT 0 685.335 0.070 685.405 ;
    RECT 0 685.475 0.070 685.545 ;
    RECT 0 685.615 0.070 685.685 ;
    RECT 0 685.755 0.070 685.825 ;
    RECT 0 685.895 0.070 685.965 ;
    RECT 0 686.035 0.070 686.105 ;
    RECT 0 686.175 0.070 686.245 ;
    RECT 0 686.315 0.070 686.385 ;
    RECT 0 686.455 0.070 686.525 ;
    RECT 0 686.595 0.070 686.665 ;
    RECT 0 686.735 0.070 686.805 ;
    RECT 0 686.875 0.070 686.945 ;
    RECT 0 687.015 0.070 687.085 ;
    RECT 0 687.155 0.070 687.225 ;
    RECT 0 687.295 0.070 687.365 ;
    RECT 0 687.435 0.070 687.505 ;
    RECT 0 687.575 0.070 687.645 ;
    RECT 0 687.715 0.070 687.785 ;
    RECT 0 687.855 0.070 687.925 ;
    RECT 0 687.995 0.070 688.065 ;
    RECT 0 688.135 0.070 688.205 ;
    RECT 0 688.275 0.070 688.345 ;
    RECT 0 688.415 0.070 688.485 ;
    RECT 0 688.555 0.070 688.625 ;
    RECT 0 688.695 0.070 688.765 ;
    RECT 0 688.835 0.070 688.905 ;
    RECT 0 688.975 0.070 689.045 ;
    RECT 0 689.115 0.070 689.185 ;
    RECT 0 689.255 0.070 689.325 ;
    RECT 0 689.395 0.070 689.465 ;
    RECT 0 689.535 0.070 689.605 ;
    RECT 0 689.675 0.070 689.745 ;
    RECT 0 689.815 0.070 689.885 ;
    RECT 0 689.955 0.070 690.025 ;
    RECT 0 690.095 0.070 690.165 ;
    RECT 0 690.235 0.070 690.305 ;
    RECT 0 690.375 0.070 690.445 ;
    RECT 0 690.515 0.070 690.585 ;
    RECT 0 690.655 0.070 690.725 ;
    RECT 0 690.795 0.070 690.865 ;
    RECT 0 690.935 0.070 691.005 ;
    RECT 0 691.075 0.070 691.145 ;
    RECT 0 691.215 0.070 691.285 ;
    RECT 0 691.355 0.070 691.425 ;
    RECT 0 691.495 0.070 691.565 ;
    RECT 0 691.635 0.070 691.705 ;
    RECT 0 691.775 0.070 691.845 ;
    RECT 0 691.915 0.070 691.985 ;
    RECT 0 692.055 0.070 692.125 ;
    RECT 0 692.195 0.070 692.265 ;
    RECT 0 692.335 0.070 692.405 ;
    RECT 0 692.475 0.070 692.545 ;
    RECT 0 692.615 0.070 692.685 ;
    RECT 0 692.755 0.070 692.825 ;
    RECT 0 692.895 0.070 692.965 ;
    RECT 0 693.035 0.070 693.105 ;
    RECT 0 693.175 0.070 693.245 ;
    RECT 0 693.315 0.070 693.385 ;
    RECT 0 693.455 0.070 693.525 ;
    RECT 0 693.595 0.070 693.665 ;
    RECT 0 693.735 0.070 693.805 ;
    RECT 0 693.875 0.070 693.945 ;
    RECT 0 694.015 0.070 694.085 ;
    RECT 0 694.155 0.070 694.225 ;
    RECT 0 694.295 0.070 694.365 ;
    RECT 0 694.435 0.070 694.505 ;
    RECT 0 694.575 0.070 694.645 ;
    RECT 0 694.715 0.070 694.785 ;
    RECT 0 694.855 0.070 694.925 ;
    RECT 0 694.995 0.070 695.065 ;
    RECT 0 695.135 0.070 695.205 ;
    RECT 0 695.275 0.070 695.345 ;
    RECT 0 695.415 0.070 695.485 ;
    RECT 0 695.555 0.070 695.625 ;
    RECT 0 695.695 0.070 695.765 ;
    RECT 0 695.835 0.070 695.905 ;
    RECT 0 695.975 0.070 696.045 ;
    RECT 0 696.115 0.070 696.185 ;
    RECT 0 696.255 0.070 696.325 ;
    RECT 0 696.395 0.070 696.465 ;
    RECT 0 696.535 0.070 696.605 ;
    RECT 0 696.675 0.070 696.745 ;
    RECT 0 696.815 0.070 696.885 ;
    RECT 0 696.955 0.070 697.025 ;
    RECT 0 697.095 0.070 697.165 ;
    RECT 0 697.235 0.070 697.305 ;
    RECT 0 697.375 0.070 697.445 ;
    RECT 0 697.515 0.070 697.585 ;
    RECT 0 697.655 0.070 697.725 ;
    RECT 0 697.795 0.070 697.865 ;
    RECT 0 697.935 0.070 698.005 ;
    RECT 0 698.075 0.070 698.145 ;
    RECT 0 698.215 0.070 698.285 ;
    RECT 0 698.355 0.070 698.425 ;
    RECT 0 698.495 0.070 698.565 ;
    RECT 0 698.635 0.070 698.705 ;
    RECT 0 698.775 0.070 698.845 ;
    RECT 0 698.915 0.070 698.985 ;
    RECT 0 699.055 0.070 699.125 ;
    RECT 0 699.195 0.070 699.265 ;
    RECT 0 699.335 0.070 699.405 ;
    RECT 0 699.475 0.070 699.545 ;
    RECT 0 699.615 0.070 699.685 ;
    RECT 0 699.755 0.070 699.825 ;
    RECT 0 699.895 0.070 699.965 ;
    RECT 0 700.035 0.070 700.105 ;
    RECT 0 700.175 0.070 700.245 ;
    RECT 0 700.315 0.070 700.385 ;
    RECT 0 700.455 0.070 700.525 ;
    RECT 0 700.595 0.070 700.665 ;
    RECT 0 700.735 0.070 700.805 ;
    RECT 0 700.875 0.070 700.945 ;
    RECT 0 701.015 0.070 701.085 ;
    RECT 0 701.155 0.070 701.225 ;
    RECT 0 701.295 0.070 701.365 ;
    RECT 0 701.435 0.070 701.505 ;
    RECT 0 701.575 0.070 701.645 ;
    RECT 0 701.715 0.070 701.785 ;
    RECT 0 701.855 0.070 701.925 ;
    RECT 0 701.995 0.070 702.065 ;
    RECT 0 702.135 0.070 702.205 ;
    RECT 0 702.275 0.070 702.345 ;
    RECT 0 702.415 0.070 702.485 ;
    RECT 0 702.555 0.070 702.625 ;
    RECT 0 702.695 0.070 702.765 ;
    RECT 0 702.835 0.070 702.905 ;
    RECT 0 702.975 0.070 703.045 ;
    RECT 0 703.115 0.070 703.185 ;
    RECT 0 703.255 0.070 703.325 ;
    RECT 0 703.395 0.070 703.465 ;
    RECT 0 703.535 0.070 703.605 ;
    RECT 0 703.675 0.070 703.745 ;
    RECT 0 703.815 0.070 703.885 ;
    RECT 0 703.955 0.070 704.025 ;
    RECT 0 704.095 0.070 704.165 ;
    RECT 0 704.235 0.070 704.305 ;
    RECT 0 704.375 0.070 704.445 ;
    RECT 0 704.515 0.070 704.585 ;
    RECT 0 704.655 0.070 704.725 ;
    RECT 0 704.795 0.070 704.865 ;
    RECT 0 704.935 0.070 705.005 ;
    RECT 0 705.075 0.070 705.145 ;
    RECT 0 705.215 0.070 705.285 ;
    RECT 0 705.355 0.070 705.425 ;
    RECT 0 705.495 0.070 705.565 ;
    RECT 0 705.635 0.070 705.705 ;
    RECT 0 705.775 0.070 705.845 ;
    RECT 0 705.915 0.070 705.985 ;
    RECT 0 706.055 0.070 706.125 ;
    RECT 0 706.195 0.070 706.265 ;
    RECT 0 706.335 0.070 706.405 ;
    RECT 0 706.475 0.070 706.545 ;
    RECT 0 706.615 0.070 706.685 ;
    RECT 0 706.755 0.070 706.825 ;
    RECT 0 706.895 0.070 706.965 ;
    RECT 0 707.035 0.070 707.105 ;
    RECT 0 707.175 0.070 707.245 ;
    RECT 0 707.315 0.070 707.385 ;
    RECT 0 707.455 0.070 707.525 ;
    RECT 0 707.595 0.070 707.665 ;
    RECT 0 707.735 0.070 707.805 ;
    RECT 0 707.875 0.070 707.945 ;
    RECT 0 708.015 0.070 708.085 ;
    RECT 0 708.155 0.070 708.225 ;
    RECT 0 708.295 0.070 708.365 ;
    RECT 0 708.435 0.070 708.505 ;
    RECT 0 708.575 0.070 708.645 ;
    RECT 0 708.715 0.070 708.785 ;
    RECT 0 708.855 0.070 708.925 ;
    RECT 0 708.995 0.070 709.065 ;
    RECT 0 709.135 0.070 709.205 ;
    RECT 0 709.275 0.070 709.345 ;
    RECT 0 709.415 0.070 709.485 ;
    RECT 0 709.555 0.070 709.625 ;
    RECT 0 709.695 0.070 709.765 ;
    RECT 0 709.835 0.070 709.905 ;
    RECT 0 709.975 0.070 710.045 ;
    RECT 0 710.115 0.070 710.185 ;
    RECT 0 710.255 0.070 710.325 ;
    RECT 0 710.395 0.070 710.465 ;
    RECT 0 710.535 0.070 710.605 ;
    RECT 0 710.675 0.070 710.745 ;
    RECT 0 710.815 0.070 710.885 ;
    RECT 0 710.955 0.070 711.025 ;
    RECT 0 711.095 0.070 711.165 ;
    RECT 0 711.235 0.070 711.305 ;
    RECT 0 711.375 0.070 711.445 ;
    RECT 0 711.515 0.070 711.585 ;
    RECT 0 711.655 0.070 711.725 ;
    RECT 0 711.795 0.070 711.865 ;
    RECT 0 711.935 0.070 712.005 ;
    RECT 0 712.075 0.070 712.145 ;
    RECT 0 712.215 0.070 712.285 ;
    RECT 0 712.355 0.070 712.425 ;
    RECT 0 712.495 0.070 712.565 ;
    RECT 0 712.635 0.070 712.705 ;
    RECT 0 712.775 0.070 712.845 ;
    RECT 0 712.915 0.070 712.985 ;
    RECT 0 713.055 0.070 713.125 ;
    RECT 0 713.195 0.070 713.265 ;
    RECT 0 713.335 0.070 713.405 ;
    RECT 0 713.475 0.070 713.545 ;
    RECT 0 713.615 0.070 713.685 ;
    RECT 0 713.755 0.070 713.825 ;
    RECT 0 713.895 0.070 713.965 ;
    RECT 0 714.035 0.070 714.105 ;
    RECT 0 714.175 0.070 714.245 ;
    RECT 0 714.315 0.070 714.385 ;
    RECT 0 714.455 0.070 714.525 ;
    RECT 0 714.595 0.070 714.665 ;
    RECT 0 714.735 0.070 714.805 ;
    RECT 0 714.875 0.070 714.945 ;
    RECT 0 715.015 0.070 715.085 ;
    RECT 0 715.155 0.070 715.225 ;
    RECT 0 715.295 0.070 715.365 ;
    RECT 0 715.435 0.070 715.505 ;
    RECT 0 715.575 0.070 715.645 ;
    RECT 0 715.715 0.070 715.785 ;
    RECT 0 715.855 0.070 715.925 ;
    RECT 0 715.995 0.070 716.065 ;
    RECT 0 716.135 0.070 716.205 ;
    RECT 0 716.275 0.070 716.345 ;
    RECT 0 716.415 0.070 716.485 ;
    RECT 0 716.555 0.070 716.625 ;
    RECT 0 716.695 0.070 716.765 ;
    RECT 0 716.835 0.070 716.905 ;
    RECT 0 716.975 0.070 717.045 ;
    RECT 0 717.115 0.070 717.185 ;
    RECT 0 717.255 0.070 717.325 ;
    RECT 0 717.395 0.070 717.465 ;
    RECT 0 717.535 0.070 717.605 ;
    RECT 0 717.675 0.070 717.745 ;
    RECT 0 717.815 0.070 717.885 ;
    RECT 0 717.955 0.070 718.025 ;
    RECT 0 718.095 0.070 718.165 ;
    RECT 0 718.235 0.070 718.305 ;
    RECT 0 718.375 0.070 718.445 ;
    RECT 0 718.515 0.070 718.585 ;
    RECT 0 718.655 0.070 718.725 ;
    RECT 0 718.795 0.070 718.865 ;
    RECT 0 718.935 0.070 719.005 ;
    RECT 0 719.075 0.070 719.145 ;
    RECT 0 719.215 0.070 719.285 ;
    RECT 0 719.355 0.070 719.425 ;
    RECT 0 719.495 0.070 719.565 ;
    RECT 0 719.635 0.070 719.705 ;
    RECT 0 719.775 0.070 719.845 ;
    RECT 0 719.915 0.070 719.985 ;
    RECT 0 720.055 0.070 720.125 ;
    RECT 0 720.195 0.070 720.265 ;
    RECT 0 720.335 0.070 720.405 ;
    RECT 0 720.475 0.070 720.545 ;
    RECT 0 720.615 0.070 720.685 ;
    RECT 0 720.755 0.070 720.825 ;
    RECT 0 720.895 0.070 720.965 ;
    RECT 0 721.035 0.070 721.105 ;
    RECT 0 721.175 0.070 721.245 ;
    RECT 0 721.315 0.070 721.385 ;
    RECT 0 721.455 0.070 721.525 ;
    RECT 0 721.595 0.070 721.665 ;
    RECT 0 721.735 0.070 721.805 ;
    RECT 0 721.875 0.070 721.945 ;
    RECT 0 722.015 0.070 722.085 ;
    RECT 0 722.155 0.070 722.225 ;
    RECT 0 722.295 0.070 722.365 ;
    RECT 0 722.435 0.070 722.505 ;
    RECT 0 722.575 0.070 722.645 ;
    RECT 0 722.715 0.070 722.785 ;
    RECT 0 722.855 0.070 722.925 ;
    RECT 0 722.995 0.070 723.065 ;
    RECT 0 723.135 0.070 723.205 ;
    RECT 0 723.275 0.070 723.345 ;
    RECT 0 723.415 0.070 723.485 ;
    RECT 0 723.555 0.070 723.625 ;
    RECT 0 723.695 0.070 723.765 ;
    RECT 0 723.835 0.070 723.905 ;
    RECT 0 723.975 0.070 724.045 ;
    RECT 0 724.115 0.070 724.185 ;
    RECT 0 724.255 0.070 724.325 ;
    RECT 0 724.395 0.070 724.465 ;
    RECT 0 724.535 0.070 724.605 ;
    RECT 0 724.675 0.070 724.745 ;
    RECT 0 724.815 0.070 724.885 ;
    RECT 0 724.955 0.070 725.025 ;
    RECT 0 725.095 0.070 725.165 ;
    RECT 0 725.235 0.070 725.305 ;
    RECT 0 725.375 0.070 725.445 ;
    RECT 0 725.515 0.070 725.585 ;
    RECT 0 725.655 0.070 725.725 ;
    RECT 0 725.795 0.070 725.865 ;
    RECT 0 725.935 0.070 726.005 ;
    RECT 0 726.075 0.070 726.145 ;
    RECT 0 726.215 0.070 726.285 ;
    RECT 0 726.355 0.070 726.425 ;
    RECT 0 726.495 0.070 726.565 ;
    RECT 0 726.635 0.070 726.705 ;
    RECT 0 726.775 0.070 726.845 ;
    RECT 0 726.915 0.070 726.985 ;
    RECT 0 727.055 0.070 727.125 ;
    RECT 0 727.195 0.070 727.265 ;
    RECT 0 727.335 0.070 727.405 ;
    RECT 0 727.475 0.070 727.545 ;
    RECT 0 727.615 0.070 727.685 ;
    RECT 0 727.755 0.070 727.825 ;
    RECT 0 727.895 0.070 727.965 ;
    RECT 0 728.035 0.070 728.105 ;
    RECT 0 728.175 0.070 728.245 ;
    RECT 0 728.315 0.070 728.385 ;
    RECT 0 728.455 0.070 728.525 ;
    RECT 0 728.595 0.070 728.665 ;
    RECT 0 728.735 0.070 728.805 ;
    RECT 0 728.875 0.070 728.945 ;
    RECT 0 729.015 0.070 729.085 ;
    RECT 0 729.155 0.070 729.225 ;
    RECT 0 729.295 0.070 729.365 ;
    RECT 0 729.435 0.070 729.505 ;
    RECT 0 729.575 0.070 729.645 ;
    RECT 0 729.715 0.070 729.785 ;
    RECT 0 729.855 0.070 729.925 ;
    RECT 0 729.995 0.070 730.065 ;
    RECT 0 730.135 0.070 730.205 ;
    RECT 0 730.275 0.070 730.345 ;
    RECT 0 730.415 0.070 730.485 ;
    RECT 0 730.555 0.070 730.625 ;
    RECT 0 730.695 0.070 730.765 ;
    RECT 0 730.835 0.070 730.905 ;
    RECT 0 730.975 0.070 731.045 ;
    RECT 0 731.115 0.070 731.185 ;
    RECT 0 731.255 0.070 731.325 ;
    RECT 0 731.395 0.070 731.465 ;
    RECT 0 731.535 0.070 731.605 ;
    RECT 0 731.675 0.070 731.745 ;
    RECT 0 731.815 0.070 731.885 ;
    RECT 0 731.955 0.070 732.025 ;
    RECT 0 732.095 0.070 732.165 ;
    RECT 0 732.235 0.070 732.305 ;
    RECT 0 732.375 0.070 732.445 ;
    RECT 0 732.515 0.070 732.585 ;
    RECT 0 732.655 0.070 732.725 ;
    RECT 0 732.795 0.070 732.865 ;
    RECT 0 732.935 0.070 733.005 ;
    RECT 0 733.075 0.070 733.145 ;
    RECT 0 733.215 0.070 733.285 ;
    RECT 0 733.355 0.070 733.425 ;
    RECT 0 733.495 0.070 733.565 ;
    RECT 0 733.635 0.070 733.705 ;
    RECT 0 733.775 0.070 733.845 ;
    RECT 0 733.915 0.070 733.985 ;
    RECT 0 734.055 0.070 734.125 ;
    RECT 0 734.195 0.070 734.265 ;
    RECT 0 734.335 0.070 734.405 ;
    RECT 0 734.475 0.070 734.545 ;
    RECT 0 734.615 0.070 734.685 ;
    RECT 0 734.755 0.070 734.825 ;
    RECT 0 734.895 0.070 734.965 ;
    RECT 0 735.035 0.070 735.105 ;
    RECT 0 735.175 0.070 735.245 ;
    RECT 0 735.315 0.070 735.385 ;
    RECT 0 735.455 0.070 735.525 ;
    RECT 0 735.595 0.070 735.665 ;
    RECT 0 735.735 0.070 735.805 ;
    RECT 0 735.875 0.070 735.945 ;
    RECT 0 736.015 0.070 736.085 ;
    RECT 0 736.155 0.070 736.225 ;
    RECT 0 736.295 0.070 736.365 ;
    RECT 0 736.435 0.070 736.505 ;
    RECT 0 736.575 0.070 736.645 ;
    RECT 0 736.715 0.070 736.785 ;
    RECT 0 736.855 0.070 736.925 ;
    RECT 0 736.995 0.070 737.065 ;
    RECT 0 737.135 0.070 737.205 ;
    RECT 0 737.275 0.070 737.345 ;
    RECT 0 737.415 0.070 737.485 ;
    RECT 0 737.555 0.070 737.625 ;
    RECT 0 737.695 0.070 737.765 ;
    RECT 0 737.835 0.070 737.905 ;
    RECT 0 737.975 0.070 738.045 ;
    RECT 0 738.115 0.070 738.185 ;
    RECT 0 738.255 0.070 738.325 ;
    RECT 0 738.395 0.070 738.465 ;
    RECT 0 738.535 0.070 738.605 ;
    RECT 0 738.675 0.070 738.745 ;
    RECT 0 738.815 0.070 738.885 ;
    RECT 0 738.955 0.070 739.025 ;
    RECT 0 739.095 0.070 739.165 ;
    RECT 0 739.235 0.070 739.305 ;
    RECT 0 739.375 0.070 739.445 ;
    RECT 0 739.515 0.070 739.585 ;
    RECT 0 739.655 0.070 739.725 ;
    RECT 0 739.795 0.070 739.865 ;
    RECT 0 739.935 0.070 740.005 ;
    RECT 0 740.075 0.070 740.145 ;
    RECT 0 740.215 0.070 740.285 ;
    RECT 0 740.355 0.070 740.425 ;
    RECT 0 740.495 0.070 740.565 ;
    RECT 0 740.635 0.070 740.705 ;
    RECT 0 740.775 0.070 740.845 ;
    RECT 0 740.915 0.070 740.985 ;
    RECT 0 741.055 0.070 741.125 ;
    RECT 0 741.195 0.070 741.265 ;
    RECT 0 741.335 0.070 741.405 ;
    RECT 0 741.475 0.070 741.545 ;
    RECT 0 741.615 0.070 741.685 ;
    RECT 0 741.755 0.070 741.825 ;
    RECT 0 741.895 0.070 741.965 ;
    RECT 0 742.035 0.070 742.105 ;
    RECT 0 742.175 0.070 742.245 ;
    RECT 0 742.315 0.070 742.385 ;
    RECT 0 742.455 0.070 742.525 ;
    RECT 0 742.595 0.070 742.665 ;
    RECT 0 742.735 0.070 742.805 ;
    RECT 0 742.875 0.070 742.945 ;
    RECT 0 743.015 0.070 743.085 ;
    RECT 0 743.155 0.070 743.225 ;
    RECT 0 743.295 0.070 743.365 ;
    RECT 0 743.435 0.070 743.505 ;
    RECT 0 743.575 0.070 743.645 ;
    RECT 0 743.715 0.070 743.785 ;
    RECT 0 743.855 0.070 743.925 ;
    RECT 0 743.995 0.070 744.065 ;
    RECT 0 744.135 0.070 744.205 ;
    RECT 0 744.275 0.070 744.345 ;
    RECT 0 744.415 0.070 744.485 ;
    RECT 0 744.555 0.070 744.625 ;
    RECT 0 744.695 0.070 744.765 ;
    RECT 0 744.835 0.070 744.905 ;
    RECT 0 744.975 0.070 745.045 ;
    RECT 0 745.115 0.070 745.185 ;
    RECT 0 745.255 0.070 745.325 ;
    RECT 0 745.395 0.070 745.465 ;
    RECT 0 745.535 0.070 745.605 ;
    RECT 0 745.675 0.070 745.745 ;
    RECT 0 745.815 0.070 745.885 ;
    RECT 0 745.955 0.070 746.025 ;
    RECT 0 746.095 0.070 746.165 ;
    RECT 0 746.235 0.070 746.305 ;
    RECT 0 746.375 0.070 746.445 ;
    RECT 0 746.515 0.070 746.585 ;
    RECT 0 746.655 0.070 746.725 ;
    RECT 0 746.795 0.070 746.865 ;
    RECT 0 746.935 0.070 747.005 ;
    RECT 0 747.075 0.070 747.145 ;
    RECT 0 747.215 0.070 747.285 ;
    RECT 0 747.355 0.070 747.425 ;
    RECT 0 747.495 0.070 747.565 ;
    RECT 0 747.635 0.070 747.705 ;
    RECT 0 747.775 0.070 747.845 ;
    RECT 0 747.915 0.070 747.985 ;
    RECT 0 748.055 0.070 748.125 ;
    RECT 0 748.195 0.070 748.265 ;
    RECT 0 748.335 0.070 748.405 ;
    RECT 0 748.475 0.070 748.545 ;
    RECT 0 748.615 0.070 748.685 ;
    RECT 0 748.755 0.070 748.825 ;
    RECT 0 748.895 0.070 748.965 ;
    RECT 0 749.035 0.070 749.105 ;
    RECT 0 749.175 0.070 749.245 ;
    RECT 0 749.315 0.070 749.385 ;
    RECT 0 749.455 0.070 749.525 ;
    RECT 0 749.595 0.070 749.665 ;
    RECT 0 749.735 0.070 749.805 ;
    RECT 0 749.875 0.070 749.945 ;
    RECT 0 750.015 0.070 750.085 ;
    RECT 0 750.155 0.070 750.225 ;
    RECT 0 750.295 0.070 750.365 ;
    RECT 0 750.435 0.070 750.505 ;
    RECT 0 750.575 0.070 750.645 ;
    RECT 0 750.715 0.070 750.785 ;
    RECT 0 750.855 0.070 750.925 ;
    RECT 0 750.995 0.070 751.065 ;
    RECT 0 751.135 0.070 751.205 ;
    RECT 0 751.275 0.070 751.345 ;
    RECT 0 751.415 0.070 751.485 ;
    RECT 0 751.555 0.070 751.625 ;
    RECT 0 751.695 0.070 751.765 ;
    RECT 0 751.835 0.070 751.905 ;
    RECT 0 751.975 0.070 752.045 ;
    RECT 0 752.115 0.070 752.185 ;
    RECT 0 752.255 0.070 752.325 ;
    RECT 0 752.395 0.070 752.465 ;
    RECT 0 752.535 0.070 752.605 ;
    RECT 0 752.675 0.070 752.745 ;
    RECT 0 752.815 0.070 752.885 ;
    RECT 0 752.955 0.070 753.025 ;
    RECT 0 753.095 0.070 753.165 ;
    RECT 0 753.235 0.070 753.305 ;
    RECT 0 753.375 0.070 753.445 ;
    RECT 0 753.515 0.070 753.585 ;
    RECT 0 753.655 0.070 753.725 ;
    RECT 0 753.795 0.070 753.865 ;
    RECT 0 753.935 0.070 754.005 ;
    RECT 0 754.075 0.070 754.145 ;
    RECT 0 754.215 0.070 754.285 ;
    RECT 0 754.355 0.070 754.425 ;
    RECT 0 754.495 0.070 754.565 ;
    RECT 0 754.635 0.070 754.705 ;
    RECT 0 754.775 0.070 754.845 ;
    RECT 0 754.915 0.070 754.985 ;
    RECT 0 755.055 0.070 755.125 ;
    RECT 0 755.195 0.070 755.265 ;
    RECT 0 755.335 0.070 755.405 ;
    RECT 0 755.475 0.070 755.545 ;
    RECT 0 755.615 0.070 755.685 ;
    RECT 0 755.755 0.070 755.825 ;
    RECT 0 755.895 0.070 755.965 ;
    RECT 0 756.035 0.070 756.105 ;
    RECT 0 756.175 0.070 756.245 ;
    RECT 0 756.315 0.070 756.385 ;
    RECT 0 756.455 0.070 756.525 ;
    RECT 0 756.595 0.070 756.665 ;
    RECT 0 756.735 0.070 756.805 ;
    RECT 0 756.875 0.070 756.945 ;
    RECT 0 757.015 0.070 757.085 ;
    RECT 0 757.155 0.070 757.225 ;
    RECT 0 757.295 0.070 757.365 ;
    RECT 0 757.435 0.070 757.505 ;
    RECT 0 757.575 0.070 757.645 ;
    RECT 0 757.715 0.070 757.785 ;
    RECT 0 757.855 0.070 757.925 ;
    RECT 0 757.995 0.070 758.065 ;
    RECT 0 758.135 0.070 758.205 ;
    RECT 0 758.275 0.070 758.345 ;
    RECT 0 758.415 0.070 758.485 ;
    RECT 0 758.555 0.070 758.625 ;
    RECT 0 758.695 0.070 758.765 ;
    RECT 0 758.835 0.070 758.905 ;
    RECT 0 758.975 0.070 759.045 ;
    RECT 0 759.115 0.070 759.185 ;
    RECT 0 759.255 0.070 759.325 ;
    RECT 0 759.395 0.070 759.465 ;
    RECT 0 759.535 0.070 759.605 ;
    RECT 0 759.675 0.070 759.745 ;
    RECT 0 759.815 0.070 759.885 ;
    RECT 0 759.955 0.070 760.025 ;
    RECT 0 760.095 0.070 760.165 ;
    RECT 0 760.235 0.070 760.305 ;
    RECT 0 760.375 0.070 760.445 ;
    RECT 0 760.515 0.070 760.585 ;
    RECT 0 760.655 0.070 760.725 ;
    RECT 0 760.795 0.070 760.865 ;
    RECT 0 760.935 0.070 761.005 ;
    RECT 0 761.075 0.070 761.145 ;
    RECT 0 761.215 0.070 761.285 ;
    RECT 0 761.355 0.070 761.425 ;
    RECT 0 761.495 0.070 761.565 ;
    RECT 0 761.635 0.070 761.705 ;
    RECT 0 761.775 0.070 761.845 ;
    RECT 0 761.915 0.070 761.985 ;
    RECT 0 762.055 0.070 762.125 ;
    RECT 0 762.195 0.070 762.265 ;
    RECT 0 762.335 0.070 762.405 ;
    RECT 0 762.475 0.070 762.545 ;
    RECT 0 762.615 0.070 762.685 ;
    RECT 0 762.755 0.070 762.825 ;
    RECT 0 762.895 0.070 762.965 ;
    RECT 0 763.035 0.070 763.105 ;
    RECT 0 763.175 0.070 763.245 ;
    RECT 0 763.315 0.070 763.385 ;
    RECT 0 763.455 0.070 763.525 ;
    RECT 0 763.595 0.070 763.665 ;
    RECT 0 763.735 0.070 763.805 ;
    RECT 0 763.875 0.070 763.945 ;
    RECT 0 764.015 0.070 764.085 ;
    RECT 0 764.155 0.070 764.225 ;
    RECT 0 764.295 0.070 764.365 ;
    RECT 0 764.435 0.070 764.505 ;
    RECT 0 764.575 0.070 764.645 ;
    RECT 0 764.715 0.070 764.785 ;
    RECT 0 764.855 0.070 764.925 ;
    RECT 0 764.995 0.070 765.065 ;
    RECT 0 765.135 0.070 765.205 ;
    RECT 0 765.275 0.070 765.345 ;
    RECT 0 765.415 0.070 765.485 ;
    RECT 0 765.555 0.070 765.625 ;
    RECT 0 765.695 0.070 765.765 ;
    RECT 0 765.835 0.070 765.905 ;
    RECT 0 765.975 0.070 766.045 ;
    RECT 0 766.115 0.070 766.185 ;
    RECT 0 766.255 0.070 766.325 ;
    RECT 0 766.395 0.070 766.465 ;
    RECT 0 766.535 0.070 766.605 ;
    RECT 0 766.675 0.070 766.745 ;
    RECT 0 766.815 0.070 766.885 ;
    RECT 0 766.955 0.070 767.025 ;
    RECT 0 767.095 0.070 767.165 ;
    RECT 0 767.235 0.070 767.305 ;
    RECT 0 767.375 0.070 767.445 ;
    RECT 0 767.515 0.070 767.585 ;
    RECT 0 767.655 0.070 767.725 ;
    RECT 0 767.795 0.070 767.865 ;
    RECT 0 767.935 0.070 768.005 ;
    RECT 0 768.075 0.070 768.145 ;
    RECT 0 768.215 0.070 768.285 ;
    RECT 0 768.355 0.070 768.425 ;
    RECT 0 768.495 0.070 768.565 ;
    RECT 0 768.635 0.070 768.705 ;
    RECT 0 768.775 0.070 768.845 ;
    RECT 0 768.915 0.070 768.985 ;
    RECT 0 769.055 0.070 769.125 ;
    RECT 0 769.195 0.070 769.265 ;
    RECT 0 769.335 0.070 769.405 ;
    RECT 0 769.475 0.070 769.545 ;
    RECT 0 769.615 0.070 769.685 ;
    RECT 0 769.755 0.070 769.825 ;
    RECT 0 769.895 0.070 769.965 ;
    RECT 0 770.035 0.070 770.105 ;
    RECT 0 770.175 0.070 770.245 ;
    RECT 0 770.315 0.070 770.385 ;
    RECT 0 770.455 0.070 770.525 ;
    RECT 0 770.595 0.070 770.665 ;
    RECT 0 770.735 0.070 770.805 ;
    RECT 0 770.875 0.070 770.945 ;
    RECT 0 771.015 0.070 771.085 ;
    RECT 0 771.155 0.070 771.225 ;
    RECT 0 771.295 0.070 771.365 ;
    RECT 0 771.435 0.070 771.505 ;
    RECT 0 771.575 0.070 771.645 ;
    RECT 0 771.715 0.070 771.785 ;
    RECT 0 771.855 0.070 771.925 ;
    RECT 0 771.995 0.070 772.065 ;
    RECT 0 772.135 0.070 772.205 ;
    RECT 0 772.275 0.070 772.345 ;
    RECT 0 772.415 0.070 772.485 ;
    RECT 0 772.555 0.070 772.625 ;
    RECT 0 772.695 0.070 772.765 ;
    RECT 0 772.835 0.070 772.905 ;
    RECT 0 772.975 0.070 773.045 ;
    RECT 0 773.115 0.070 773.185 ;
    RECT 0 773.255 0.070 773.325 ;
    RECT 0 773.395 0.070 773.465 ;
    RECT 0 773.535 0.070 773.605 ;
    RECT 0 773.675 0.070 773.745 ;
    RECT 0 773.815 0.070 773.885 ;
    RECT 0 773.955 0.070 774.025 ;
    RECT 0 774.095 0.070 774.165 ;
    RECT 0 774.235 0.070 774.305 ;
    RECT 0 774.375 0.070 774.445 ;
    RECT 0 774.515 0.070 774.585 ;
    RECT 0 774.655 0.070 774.725 ;
    RECT 0 774.795 0.070 774.865 ;
    RECT 0 774.935 0.070 775.005 ;
    RECT 0 775.075 0.070 775.145 ;
    RECT 0 775.215 0.070 775.285 ;
    RECT 0 775.355 0.070 775.425 ;
    RECT 0 775.495 0.070 775.565 ;
    RECT 0 775.635 0.070 775.705 ;
    RECT 0 775.775 0.070 775.845 ;
    RECT 0 775.915 0.070 775.985 ;
    RECT 0 776.055 0.070 776.125 ;
    RECT 0 776.195 0.070 776.265 ;
    RECT 0 776.335 0.070 776.405 ;
    RECT 0 776.475 0.070 776.545 ;
    RECT 0 776.615 0.070 776.685 ;
    RECT 0 776.755 0.070 776.825 ;
    RECT 0 776.895 0.070 776.965 ;
    RECT 0 777.035 0.070 777.105 ;
    RECT 0 777.175 0.070 777.245 ;
    RECT 0 777.315 0.070 777.385 ;
    RECT 0 777.455 0.070 777.525 ;
    RECT 0 777.595 0.070 777.665 ;
    RECT 0 777.735 0.070 777.805 ;
    RECT 0 777.875 0.070 777.945 ;
    RECT 0 778.015 0.070 778.085 ;
    RECT 0 778.155 0.070 778.225 ;
    RECT 0 778.295 0.070 778.365 ;
    RECT 0 778.435 0.070 778.505 ;
    RECT 0 778.575 0.070 778.645 ;
    RECT 0 778.715 0.070 778.785 ;
    RECT 0 778.855 0.070 778.925 ;
    RECT 0 778.995 0.070 779.065 ;
    RECT 0 779.135 0.070 779.205 ;
    RECT 0 779.275 0.070 779.345 ;
    RECT 0 779.415 0.070 779.485 ;
    RECT 0 779.555 0.070 779.625 ;
    RECT 0 779.695 0.070 779.765 ;
    RECT 0 779.835 0.070 779.905 ;
    RECT 0 779.975 0.070 780.045 ;
    RECT 0 780.115 0.070 780.185 ;
    RECT 0 780.255 0.070 780.325 ;
    RECT 0 780.395 0.070 780.465 ;
    RECT 0 780.535 0.070 780.605 ;
    RECT 0 780.675 0.070 780.745 ;
    RECT 0 780.815 0.070 780.885 ;
    RECT 0 780.955 0.070 781.025 ;
    RECT 0 781.095 0.070 781.165 ;
    RECT 0 781.235 0.070 781.305 ;
    RECT 0 781.375 0.070 781.445 ;
    RECT 0 781.515 0.070 781.585 ;
    RECT 0 781.655 0.070 781.725 ;
    RECT 0 781.795 0.070 781.865 ;
    RECT 0 781.935 0.070 782.005 ;
    RECT 0 782.075 0.070 782.145 ;
    RECT 0 782.215 0.070 782.285 ;
    RECT 0 782.355 0.070 782.425 ;
    RECT 0 782.495 0.070 782.565 ;
    RECT 0 782.635 0.070 782.705 ;
    RECT 0 782.775 0.070 782.845 ;
    RECT 0 782.915 0.070 782.985 ;
    RECT 0 783.055 0.070 783.125 ;
    RECT 0 783.195 0.070 783.265 ;
    RECT 0 783.335 0.070 783.405 ;
    RECT 0 783.475 0.070 783.545 ;
    RECT 0 783.615 0.070 783.685 ;
    RECT 0 783.755 0.070 783.825 ;
    RECT 0 783.895 0.070 783.965 ;
    RECT 0 784.035 0.070 784.105 ;
    RECT 0 784.175 0.070 784.245 ;
    RECT 0 784.315 0.070 784.385 ;
    RECT 0 784.455 0.070 784.525 ;
    RECT 0 784.595 0.070 784.665 ;
    RECT 0 784.735 0.070 784.805 ;
    RECT 0 784.875 0.070 784.945 ;
    RECT 0 785.015 0.070 785.085 ;
    RECT 0 785.155 0.070 785.225 ;
    RECT 0 785.295 0.070 785.365 ;
    RECT 0 785.435 0.070 785.505 ;
    RECT 0 785.575 0.070 785.645 ;
    RECT 0 785.715 0.070 785.785 ;
    RECT 0 785.855 0.070 785.925 ;
    RECT 0 785.995 0.070 786.065 ;
    RECT 0 786.135 0.070 786.205 ;
    RECT 0 786.275 0.070 786.345 ;
    RECT 0 786.415 0.070 786.485 ;
    RECT 0 786.555 0.070 786.625 ;
    RECT 0 786.695 0.070 786.765 ;
    RECT 0 786.835 0.070 786.905 ;
    RECT 0 786.975 0.070 787.045 ;
    RECT 0 787.115 0.070 787.185 ;
    RECT 0 787.255 0.070 787.325 ;
    RECT 0 787.395 0.070 787.465 ;
    RECT 0 787.535 0.070 787.605 ;
    RECT 0 787.675 0.070 787.745 ;
    RECT 0 787.815 0.070 787.885 ;
    RECT 0 787.955 0.070 788.025 ;
    RECT 0 788.095 0.070 788.165 ;
    RECT 0 788.235 0.070 788.305 ;
    RECT 0 788.375 0.070 788.445 ;
    RECT 0 788.515 0.070 788.585 ;
    RECT 0 788.655 0.070 788.725 ;
    RECT 0 788.795 0.070 788.865 ;
    RECT 0 788.935 0.070 789.005 ;
    RECT 0 789.075 0.070 789.145 ;
    RECT 0 789.215 0.070 789.285 ;
    RECT 0 789.355 0.070 789.425 ;
    RECT 0 789.495 0.070 789.565 ;
    RECT 0 789.635 0.070 789.705 ;
    RECT 0 789.775 0.070 789.845 ;
    RECT 0 789.915 0.070 789.985 ;
    RECT 0 790.055 0.070 790.125 ;
    RECT 0 790.195 0.070 790.265 ;
    RECT 0 790.335 0.070 790.405 ;
    RECT 0 790.475 0.070 790.545 ;
    RECT 0 790.615 0.070 790.685 ;
    RECT 0 790.755 0.070 790.825 ;
    RECT 0 790.895 0.070 790.965 ;
    RECT 0 791.035 0.070 791.105 ;
    RECT 0 791.175 0.070 791.245 ;
    RECT 0 791.315 0.070 791.385 ;
    RECT 0 791.455 0.070 791.525 ;
    RECT 0 791.595 0.070 791.665 ;
    RECT 0 791.735 0.070 791.805 ;
    RECT 0 791.875 0.070 791.945 ;
    RECT 0 792.015 0.070 792.085 ;
    RECT 0 792.155 0.070 792.225 ;
    RECT 0 792.295 0.070 792.365 ;
    RECT 0 792.435 0.070 792.505 ;
    RECT 0 792.575 0.070 792.645 ;
    RECT 0 792.715 0.070 792.785 ;
    RECT 0 792.855 0.070 792.925 ;
    RECT 0 792.995 0.070 793.065 ;
    RECT 0 793.135 0.070 793.205 ;
    RECT 0 793.275 0.070 793.345 ;
    RECT 0 793.415 0.070 793.485 ;
    RECT 0 793.555 0.070 793.625 ;
    RECT 0 793.695 0.070 793.765 ;
    RECT 0 793.835 0.070 793.905 ;
    RECT 0 793.975 0.070 794.045 ;
    RECT 0 794.115 0.070 794.185 ;
    RECT 0 794.255 0.070 794.325 ;
    RECT 0 794.395 0.070 794.465 ;
    RECT 0 794.535 0.070 794.605 ;
    RECT 0 794.675 0.070 794.745 ;
    RECT 0 794.815 0.070 794.885 ;
    RECT 0 794.955 0.070 795.025 ;
    RECT 0 795.095 0.070 795.165 ;
    RECT 0 795.235 0.070 795.305 ;
    RECT 0 795.375 0.070 795.445 ;
    RECT 0 795.515 0.070 795.585 ;
    RECT 0 795.655 0.070 795.725 ;
    RECT 0 795.795 0.070 795.865 ;
    RECT 0 795.935 0.070 796.005 ;
    RECT 0 796.075 0.070 796.145 ;
    RECT 0 796.215 0.070 796.285 ;
    RECT 0 796.355 0.070 796.425 ;
    RECT 0 796.495 0.070 796.565 ;
    RECT 0 796.635 0.070 796.705 ;
    RECT 0 796.775 0.070 796.845 ;
    RECT 0 796.915 0.070 796.985 ;
    RECT 0 797.055 0.070 797.125 ;
    RECT 0 797.195 0.070 797.265 ;
    RECT 0 797.335 0.070 797.405 ;
    RECT 0 797.475 0.070 797.545 ;
    RECT 0 797.615 0.070 797.685 ;
    RECT 0 797.755 0.070 797.825 ;
    RECT 0 797.895 0.070 797.965 ;
    RECT 0 798.035 0.070 798.105 ;
    RECT 0 798.175 0.070 798.245 ;
    RECT 0 798.315 0.070 798.385 ;
    RECT 0 798.455 0.070 798.525 ;
    RECT 0 798.595 0.070 798.665 ;
    RECT 0 798.735 0.070 798.805 ;
    RECT 0 798.875 0.070 798.945 ;
    RECT 0 799.015 0.070 799.085 ;
    RECT 0 799.155 0.070 799.225 ;
    RECT 0 799.295 0.070 799.365 ;
    RECT 0 799.435 0.070 799.505 ;
    RECT 0 799.575 0.070 799.645 ;
    RECT 0 799.715 0.070 799.785 ;
    RECT 0 799.855 0.070 799.925 ;
    RECT 0 799.995 0.070 800.065 ;
    RECT 0 800.135 0.070 800.205 ;
    RECT 0 800.275 0.070 800.345 ;
    RECT 0 800.415 0.070 800.485 ;
    RECT 0 800.555 0.070 800.625 ;
    RECT 0 800.695 0.070 800.765 ;
    RECT 0 800.835 0.070 800.905 ;
    RECT 0 800.975 0.070 801.045 ;
    RECT 0 801.115 0.070 801.185 ;
    RECT 0 801.255 0.070 801.325 ;
    RECT 0 801.395 0.070 801.465 ;
    RECT 0 801.535 0.070 801.605 ;
    RECT 0 801.675 0.070 801.745 ;
    RECT 0 801.815 0.070 801.885 ;
    RECT 0 801.955 0.070 802.025 ;
    RECT 0 802.095 0.070 802.165 ;
    RECT 0 802.235 0.070 802.305 ;
    RECT 0 802.375 0.070 802.445 ;
    RECT 0 802.515 0.070 802.585 ;
    RECT 0 802.655 0.070 802.725 ;
    RECT 0 802.795 0.070 802.865 ;
    RECT 0 802.935 0.070 803.005 ;
    RECT 0 803.075 0.070 803.145 ;
    RECT 0 803.215 0.070 803.285 ;
    RECT 0 803.355 0.070 803.425 ;
    RECT 0 803.495 0.070 803.565 ;
    RECT 0 803.635 0.070 803.705 ;
    RECT 0 803.775 0.070 803.845 ;
    RECT 0 803.915 0.070 803.985 ;
    RECT 0 804.055 0.070 804.125 ;
    RECT 0 804.195 0.070 804.265 ;
    RECT 0 804.335 0.070 804.405 ;
    RECT 0 804.475 0.070 804.545 ;
    RECT 0 804.615 0.070 804.685 ;
    RECT 0 804.755 0.070 804.825 ;
    RECT 0 804.895 0.070 804.965 ;
    RECT 0 805.035 0.070 805.105 ;
    RECT 0 805.175 0.070 805.245 ;
    RECT 0 805.315 0.070 805.385 ;
    RECT 0 805.455 0.070 805.525 ;
    RECT 0 805.595 0.070 805.665 ;
    RECT 0 805.735 0.070 805.805 ;
    RECT 0 805.875 0.070 805.945 ;
    RECT 0 806.015 0.070 806.085 ;
    RECT 0 806.155 0.070 806.225 ;
    RECT 0 806.295 0.070 806.365 ;
    RECT 0 806.435 0.070 806.505 ;
    RECT 0 806.575 0.070 806.645 ;
    RECT 0 806.715 0.070 806.785 ;
    RECT 0 806.855 0.070 806.925 ;
    RECT 0 806.995 0.070 807.065 ;
    RECT 0 807.135 0.070 807.205 ;
    RECT 0 807.275 0.070 807.345 ;
    RECT 0 807.415 0.070 807.485 ;
    RECT 0 807.555 0.070 807.625 ;
    RECT 0 807.695 0.070 807.765 ;
    RECT 0 807.835 0.070 807.905 ;
    RECT 0 807.975 0.070 808.045 ;
    RECT 0 808.115 0.070 808.185 ;
    RECT 0 808.255 0.070 808.325 ;
    RECT 0 808.395 0.070 808.465 ;
    RECT 0 808.535 0.070 808.605 ;
    RECT 0 808.675 0.070 808.745 ;
    RECT 0 808.815 0.070 808.885 ;
    RECT 0 808.955 0.070 809.025 ;
    RECT 0 809.095 0.070 809.165 ;
    RECT 0 809.235 0.070 809.305 ;
    RECT 0 809.375 0.070 809.445 ;
    RECT 0 809.515 0.070 809.585 ;
    RECT 0 809.655 0.070 809.725 ;
    RECT 0 809.795 0.070 809.865 ;
    RECT 0 809.935 0.070 810.005 ;
    RECT 0 810.075 0.070 810.145 ;
    RECT 0 810.215 0.070 810.285 ;
    RECT 0 810.355 0.070 810.425 ;
    RECT 0 810.495 0.070 810.565 ;
    RECT 0 810.635 0.070 810.705 ;
    RECT 0 810.775 0.070 810.845 ;
    RECT 0 810.915 0.070 810.985 ;
    RECT 0 811.055 0.070 811.125 ;
    RECT 0 811.195 0.070 811.265 ;
    RECT 0 811.335 0.070 811.405 ;
    RECT 0 811.475 0.070 811.545 ;
    RECT 0 811.615 0.070 811.685 ;
    RECT 0 811.755 0.070 811.825 ;
    RECT 0 811.895 0.070 811.965 ;
    RECT 0 812.035 0.070 812.105 ;
    RECT 0 812.175 0.070 812.245 ;
    RECT 0 812.315 0.070 812.385 ;
    RECT 0 812.455 0.070 812.525 ;
    RECT 0 812.595 0.070 812.665 ;
    RECT 0 812.735 0.070 812.805 ;
    RECT 0 812.875 0.070 812.945 ;
    RECT 0 813.015 0.070 813.085 ;
    RECT 0 813.155 0.070 813.225 ;
    RECT 0 813.295 0.070 813.365 ;
    RECT 0 813.435 0.070 813.505 ;
    RECT 0 813.575 0.070 813.645 ;
    RECT 0 813.715 0.070 813.785 ;
    RECT 0 813.855 0.070 813.925 ;
    RECT 0 813.995 0.070 814.065 ;
    RECT 0 814.135 0.070 814.205 ;
    RECT 0 814.275 0.070 814.345 ;
    RECT 0 814.415 0.070 814.485 ;
    RECT 0 814.555 0.070 814.625 ;
    RECT 0 814.695 0.070 814.765 ;
    RECT 0 814.835 0.070 814.905 ;
    RECT 0 814.975 0.070 815.045 ;
    RECT 0 815.115 0.070 815.185 ;
    RECT 0 815.255 0.070 815.325 ;
    RECT 0 815.395 0.070 815.465 ;
    RECT 0 815.535 0.070 815.605 ;
    RECT 0 815.675 0.070 815.745 ;
    RECT 0 815.815 0.070 815.885 ;
    RECT 0 815.955 0.070 816.025 ;
    RECT 0 816.095 0.070 816.165 ;
    RECT 0 816.235 0.070 816.305 ;
    RECT 0 816.375 0.070 816.445 ;
    RECT 0 816.515 0.070 816.585 ;
    RECT 0 816.655 0.070 816.725 ;
    RECT 0 816.795 0.070 816.865 ;
    RECT 0 816.935 0.070 817.005 ;
    RECT 0 817.075 0.070 817.145 ;
    RECT 0 817.215 0.070 817.285 ;
    RECT 0 817.355 0.070 817.425 ;
    RECT 0 817.495 0.070 817.565 ;
    RECT 0 817.635 0.070 817.705 ;
    RECT 0 817.775 0.070 817.845 ;
    RECT 0 817.915 0.070 817.985 ;
    RECT 0 818.055 0.070 818.125 ;
    RECT 0 818.195 0.070 818.265 ;
    RECT 0 818.335 0.070 818.405 ;
    RECT 0 818.475 0.070 818.545 ;
    RECT 0 818.615 0.070 818.685 ;
    RECT 0 818.755 0.070 818.825 ;
    RECT 0 818.895 0.070 818.965 ;
    RECT 0 819.035 0.070 819.105 ;
    RECT 0 819.175 0.070 819.245 ;
    RECT 0 819.315 0.070 819.385 ;
    RECT 0 819.455 0.070 819.525 ;
    RECT 0 819.595 0.070 819.665 ;
    RECT 0 819.735 0.070 819.805 ;
    RECT 0 819.875 0.070 819.945 ;
    RECT 0 820.015 0.070 820.085 ;
    RECT 0 820.155 0.070 820.225 ;
    RECT 0 820.295 0.070 820.365 ;
    RECT 0 820.435 0.070 820.505 ;
    RECT 0 820.575 0.070 820.645 ;
    RECT 0 820.715 0.070 820.785 ;
    RECT 0 820.855 0.070 820.925 ;
    RECT 0 820.995 0.070 821.065 ;
    RECT 0 821.135 0.070 821.205 ;
    RECT 0 821.275 0.070 821.345 ;
    RECT 0 821.415 0.070 821.485 ;
    RECT 0 821.555 0.070 821.625 ;
    RECT 0 821.695 0.070 821.765 ;
    RECT 0 821.835 0.070 821.905 ;
    RECT 0 821.975 0.070 822.045 ;
    RECT 0 822.115 0.070 822.185 ;
    RECT 0 822.255 0.070 822.325 ;
    RECT 0 822.395 0.070 822.465 ;
    RECT 0 822.535 0.070 822.605 ;
    RECT 0 822.675 0.070 822.745 ;
    RECT 0 822.815 0.070 822.885 ;
    RECT 0 822.955 0.070 823.025 ;
    RECT 0 823.095 0.070 823.165 ;
    RECT 0 823.235 0.070 823.305 ;
    RECT 0 823.375 0.070 823.445 ;
    RECT 0 823.515 0.070 823.585 ;
    RECT 0 823.655 0.070 823.725 ;
    RECT 0 823.795 0.070 823.865 ;
    RECT 0 823.935 0.070 824.005 ;
    RECT 0 824.075 0.070 824.145 ;
    RECT 0 824.215 0.070 824.285 ;
    RECT 0 824.355 0.070 824.425 ;
    RECT 0 824.495 0.070 824.565 ;
    RECT 0 824.635 0.070 824.705 ;
    RECT 0 824.775 0.070 824.845 ;
    RECT 0 824.915 0.070 824.985 ;
    RECT 0 825.055 0.070 825.125 ;
    RECT 0 825.195 0.070 825.265 ;
    RECT 0 825.335 0.070 825.405 ;
    RECT 0 825.475 0.070 825.545 ;
    RECT 0 825.615 0.070 825.685 ;
    RECT 0 825.755 0.070 825.825 ;
    RECT 0 825.895 0.070 825.965 ;
    RECT 0 826.035 0.070 826.105 ;
    RECT 0 826.175 0.070 826.245 ;
    RECT 0 826.315 0.070 826.385 ;
    RECT 0 826.455 0.070 826.525 ;
    RECT 0 826.595 0.070 826.665 ;
    RECT 0 826.735 0.070 826.805 ;
    RECT 0 826.875 0.070 826.945 ;
    RECT 0 827.015 0.070 827.085 ;
    RECT 0 827.155 0.070 827.225 ;
    RECT 0 827.295 0.070 827.365 ;
    RECT 0 827.435 0.070 827.505 ;
    RECT 0 827.575 0.070 827.645 ;
    RECT 0 827.715 0.070 827.785 ;
    RECT 0 827.855 0.070 827.925 ;
    RECT 0 827.995 0.070 828.065 ;
    RECT 0 828.135 0.070 828.205 ;
    RECT 0 828.275 0.070 828.345 ;
    RECT 0 828.415 0.070 828.485 ;
    RECT 0 828.555 0.070 828.625 ;
    RECT 0 828.695 0.070 828.765 ;
    RECT 0 828.835 0.070 828.905 ;
    RECT 0 828.975 0.070 829.045 ;
    RECT 0 829.115 0.070 829.185 ;
    RECT 0 829.255 0.070 829.325 ;
    RECT 0 829.395 0.070 829.465 ;
    RECT 0 829.535 0.070 829.605 ;
    RECT 0 829.675 0.070 829.745 ;
    RECT 0 829.815 0.070 829.885 ;
    RECT 0 829.955 0.070 830.025 ;
    RECT 0 830.095 0.070 830.165 ;
    RECT 0 830.235 0.070 830.305 ;
    RECT 0 830.375 0.070 830.445 ;
    RECT 0 830.515 0.070 830.585 ;
    RECT 0 830.655 0.070 830.725 ;
    RECT 0 830.795 0.070 830.865 ;
    RECT 0 830.935 0.070 831.005 ;
    RECT 0 831.075 0.070 831.145 ;
    RECT 0 831.215 0.070 831.285 ;
    RECT 0 831.355 0.070 831.425 ;
    RECT 0 831.495 0.070 831.565 ;
    RECT 0 831.635 0.070 831.705 ;
    RECT 0 831.775 0.070 831.845 ;
    RECT 0 831.915 0.070 831.985 ;
    RECT 0 832.055 0.070 832.125 ;
    RECT 0 832.195 0.070 832.265 ;
    RECT 0 832.335 0.070 832.405 ;
    RECT 0 832.475 0.070 832.545 ;
    RECT 0 832.615 0.070 832.685 ;
    RECT 0 832.755 0.070 832.825 ;
    RECT 0 832.895 0.070 832.965 ;
    RECT 0 833.035 0.070 833.105 ;
    RECT 0 833.175 0.070 833.245 ;
    RECT 0 833.315 0.070 833.385 ;
    RECT 0 833.455 0.070 833.525 ;
    RECT 0 833.595 0.070 833.665 ;
    RECT 0 833.735 0.070 833.805 ;
    RECT 0 833.875 0.070 833.945 ;
    RECT 0 834.015 0.070 834.085 ;
    RECT 0 834.155 0.070 834.225 ;
    RECT 0 834.295 0.070 834.365 ;
    RECT 0 834.435 0.070 834.505 ;
    RECT 0 834.575 0.070 834.645 ;
    RECT 0 834.715 0.070 834.785 ;
    RECT 0 834.855 0.070 834.925 ;
    RECT 0 834.995 0.070 835.065 ;
    RECT 0 835.135 0.070 835.205 ;
    RECT 0 835.275 0.070 835.345 ;
    RECT 0 835.415 0.070 835.485 ;
    RECT 0 835.555 0.070 835.625 ;
    RECT 0 835.695 0.070 835.765 ;
    RECT 0 835.835 0.070 835.905 ;
    RECT 0 835.975 0.070 836.045 ;
    RECT 0 836.115 0.070 836.185 ;
    RECT 0 836.255 0.070 836.325 ;
    RECT 0 836.395 0.070 836.465 ;
    RECT 0 836.535 0.070 836.605 ;
    RECT 0 836.675 0.070 836.745 ;
    RECT 0 836.815 0.070 836.885 ;
    RECT 0 836.955 0.070 837.025 ;
    RECT 0 837.095 0.070 837.165 ;
    RECT 0 837.235 0.070 837.305 ;
    RECT 0 837.375 0.070 837.445 ;
    RECT 0 837.515 0.070 837.585 ;
    RECT 0 837.655 0.070 837.725 ;
    RECT 0 837.795 0.070 837.865 ;
    RECT 0 837.935 0.070 838.005 ;
    RECT 0 838.075 0.070 838.145 ;
    RECT 0 838.215 0.070 838.285 ;
    RECT 0 838.355 0.070 838.425 ;
    RECT 0 838.495 0.070 838.565 ;
    RECT 0 838.635 0.070 838.705 ;
    RECT 0 838.775 0.070 838.845 ;
    RECT 0 838.915 0.070 838.985 ;
    RECT 0 839.055 0.070 839.125 ;
    RECT 0 839.195 0.070 839.265 ;
    RECT 0 839.335 0.070 839.405 ;
    RECT 0 839.475 0.070 839.545 ;
    RECT 0 839.615 0.070 839.685 ;
    RECT 0 839.755 0.070 839.825 ;
    RECT 0 839.895 0.070 839.965 ;
    RECT 0 840.035 0.070 840.105 ;
    RECT 0 840.175 0.070 840.245 ;
    RECT 0 840.315 0.070 840.385 ;
    RECT 0 840.455 0.070 840.525 ;
    RECT 0 840.595 0.070 840.665 ;
    RECT 0 840.735 0.070 840.805 ;
    RECT 0 840.875 0.070 840.945 ;
    RECT 0 841.015 0.070 841.085 ;
    RECT 0 841.155 0.070 841.225 ;
    RECT 0 841.295 0.070 841.365 ;
    RECT 0 841.435 0.070 841.505 ;
    RECT 0 841.575 0.070 841.645 ;
    RECT 0 841.715 0.070 841.785 ;
    RECT 0 841.855 0.070 841.925 ;
    RECT 0 841.995 0.070 842.065 ;
    RECT 0 842.135 0.070 842.205 ;
    RECT 0 842.275 0.070 842.345 ;
    RECT 0 842.415 0.070 842.485 ;
    RECT 0 842.555 0.070 842.625 ;
    RECT 0 842.695 0.070 842.765 ;
    RECT 0 842.835 0.070 842.905 ;
    RECT 0 842.975 0.070 843.045 ;
    RECT 0 843.115 0.070 843.185 ;
    RECT 0 843.255 0.070 843.325 ;
    RECT 0 843.395 0.070 843.465 ;
    RECT 0 843.535 0.070 843.605 ;
    RECT 0 843.675 0.070 843.745 ;
    RECT 0 843.815 0.070 843.885 ;
    RECT 0 843.955 0.070 844.025 ;
    RECT 0 844.095 0.070 844.165 ;
    RECT 0 844.235 0.070 844.305 ;
    RECT 0 844.375 0.070 844.445 ;
    RECT 0 844.515 0.070 844.585 ;
    RECT 0 844.655 0.070 844.725 ;
    RECT 0 844.795 0.070 844.865 ;
    RECT 0 844.935 0.070 845.005 ;
    RECT 0 845.075 0.070 845.145 ;
    RECT 0 845.215 0.070 845.285 ;
    RECT 0 845.355 0.070 845.425 ;
    RECT 0 845.495 0.070 845.565 ;
    RECT 0 845.635 0.070 845.705 ;
    RECT 0 845.775 0.070 845.845 ;
    RECT 0 845.915 0.070 845.985 ;
    RECT 0 846.055 0.070 846.125 ;
    RECT 0 846.195 0.070 846.265 ;
    RECT 0 846.335 0.070 846.405 ;
    RECT 0 846.475 0.070 846.545 ;
    RECT 0 846.615 0.070 846.685 ;
    RECT 0 846.755 0.070 846.825 ;
    RECT 0 846.895 0.070 846.965 ;
    RECT 0 847.035 0.070 847.105 ;
    RECT 0 847.175 0.070 847.245 ;
    RECT 0 847.315 0.070 847.385 ;
    RECT 0 847.455 0.070 847.525 ;
    RECT 0 847.595 0.070 847.665 ;
    RECT 0 847.735 0.070 847.805 ;
    RECT 0 847.875 0.070 847.945 ;
    RECT 0 848.015 0.070 848.085 ;
    RECT 0 848.155 0.070 848.225 ;
    RECT 0 848.295 0.070 848.365 ;
    RECT 0 848.435 0.070 848.505 ;
    RECT 0 848.575 0.070 848.645 ;
    RECT 0 848.715 0.070 848.785 ;
    RECT 0 848.855 0.070 848.925 ;
    RECT 0 848.995 0.070 849.065 ;
    RECT 0 849.135 0.070 849.205 ;
    RECT 0 849.275 0.070 849.345 ;
    RECT 0 849.415 0.070 849.485 ;
    RECT 0 849.555 0.070 849.625 ;
    RECT 0 849.695 0.070 849.765 ;
    RECT 0 849.835 0.070 849.905 ;
    RECT 0 849.975 0.070 850.045 ;
    RECT 0 850.115 0.070 850.185 ;
    RECT 0 850.255 0.070 850.325 ;
    RECT 0 850.395 0.070 850.465 ;
    RECT 0 850.535 0.070 850.605 ;
    RECT 0 850.675 0.070 850.745 ;
    RECT 0 850.815 0.070 850.885 ;
    RECT 0 850.955 0.070 851.025 ;
    RECT 0 851.095 0.070 851.165 ;
    RECT 0 851.235 0.070 851.305 ;
    RECT 0 851.375 0.070 851.445 ;
    RECT 0 851.515 0.070 851.585 ;
    RECT 0 851.655 0.070 851.725 ;
    RECT 0 851.795 0.070 851.865 ;
    RECT 0 851.935 0.070 852.005 ;
    RECT 0 852.075 0.070 852.145 ;
    RECT 0 852.215 0.070 852.285 ;
    RECT 0 852.355 0.070 852.425 ;
    RECT 0 852.495 0.070 852.565 ;
    RECT 0 852.635 0.070 852.705 ;
    RECT 0 852.775 0.070 852.845 ;
    RECT 0 852.915 0.070 852.985 ;
    RECT 0 853.055 0.070 853.125 ;
    RECT 0 853.195 0.070 853.265 ;
    RECT 0 853.335 0.070 853.405 ;
    RECT 0 853.475 0.070 853.545 ;
    RECT 0 853.615 0.070 853.685 ;
    RECT 0 853.755 0.070 853.825 ;
    RECT 0 853.895 0.070 853.965 ;
    RECT 0 854.035 0.070 854.105 ;
    RECT 0 854.175 0.070 854.245 ;
    RECT 0 854.315 0.070 854.385 ;
    RECT 0 854.455 0.070 854.525 ;
    RECT 0 854.595 0.070 854.665 ;
    RECT 0 854.735 0.070 854.805 ;
    RECT 0 854.875 0.070 854.945 ;
    RECT 0 855.015 0.070 855.085 ;
    RECT 0 855.155 0.070 855.225 ;
    RECT 0 855.295 0.070 855.365 ;
    RECT 0 855.435 0.070 855.505 ;
    RECT 0 855.575 0.070 855.645 ;
    RECT 0 855.715 0.070 855.785 ;
    RECT 0 855.855 0.070 855.925 ;
    RECT 0 855.995 0.070 856.065 ;
    RECT 0 856.135 0.070 856.205 ;
    RECT 0 856.275 0.070 856.345 ;
    RECT 0 856.415 0.070 856.485 ;
    RECT 0 856.555 0.070 856.625 ;
    RECT 0 856.695 0.070 856.765 ;
    RECT 0 856.835 0.070 856.905 ;
    RECT 0 856.975 0.070 857.045 ;
    RECT 0 857.115 0.070 857.185 ;
    RECT 0 857.255 0.070 857.325 ;
    RECT 0 857.395 0.070 857.465 ;
    RECT 0 857.535 0.070 857.605 ;
    RECT 0 857.675 0.070 857.745 ;
    RECT 0 857.815 0.070 857.885 ;
    RECT 0 857.955 0.070 858.025 ;
    RECT 0 858.095 0.070 858.165 ;
    RECT 0 858.235 0.070 858.305 ;
    RECT 0 858.375 0.070 858.445 ;
    RECT 0 858.515 0.070 858.585 ;
    RECT 0 858.655 0.070 858.725 ;
    RECT 0 858.795 0.070 858.865 ;
    RECT 0 858.935 0.070 859.005 ;
    RECT 0 859.075 0.070 859.145 ;
    RECT 0 859.215 0.070 859.285 ;
    RECT 0 859.355 0.070 859.425 ;
    RECT 0 859.495 0.070 859.565 ;
    RECT 0 859.635 0.070 859.705 ;
    RECT 0 859.775 0.070 859.845 ;
    RECT 0 859.915 0.070 859.985 ;
    RECT 0 860.055 0.070 860.125 ;
    RECT 0 860.195 0.070 860.265 ;
    RECT 0 860.335 0.070 860.405 ;
    RECT 0 860.475 0.070 860.545 ;
    RECT 0 860.615 0.070 860.685 ;
    RECT 0 860.755 0.070 860.825 ;
    RECT 0 860.895 0.070 860.965 ;
    RECT 0 861.035 0.070 861.105 ;
    RECT 0 861.175 0.070 861.245 ;
    RECT 0 861.315 0.070 861.385 ;
    RECT 0 861.455 0.070 861.525 ;
    RECT 0 861.595 0.070 861.665 ;
    RECT 0 861.735 0.070 861.805 ;
    RECT 0 861.875 0.070 861.945 ;
    RECT 0 862.015 0.070 862.085 ;
    RECT 0 862.155 0.070 862.225 ;
    RECT 0 862.295 0.070 862.365 ;
    RECT 0 862.435 0.070 862.505 ;
    RECT 0 862.575 0.070 862.645 ;
    RECT 0 862.715 0.070 862.785 ;
    RECT 0 862.855 0.070 862.925 ;
    RECT 0 862.995 0.070 863.065 ;
    RECT 0 863.135 0.070 863.205 ;
    RECT 0 863.275 0.070 863.345 ;
    RECT 0 863.415 0.070 863.485 ;
    RECT 0 863.555 0.070 863.625 ;
    RECT 0 863.695 0.070 863.765 ;
    RECT 0 863.835 0.070 863.905 ;
    RECT 0 863.975 0.070 864.045 ;
    RECT 0 864.115 0.070 864.185 ;
    RECT 0 864.255 0.070 864.325 ;
    RECT 0 864.395 0.070 864.465 ;
    RECT 0 864.535 0.070 864.605 ;
    RECT 0 864.675 0.070 864.745 ;
    RECT 0 864.815 0.070 864.885 ;
    RECT 0 864.955 0.070 865.025 ;
    RECT 0 865.095 0.070 865.165 ;
    RECT 0 865.235 0.070 865.305 ;
    RECT 0 865.375 0.070 865.445 ;
    RECT 0 865.515 0.070 865.585 ;
    RECT 0 865.655 0.070 865.725 ;
    RECT 0 865.795 0.070 865.865 ;
    RECT 0 865.935 0.070 866.005 ;
    RECT 0 866.075 0.070 866.145 ;
    RECT 0 866.215 0.070 866.285 ;
    RECT 0 866.355 0.070 866.425 ;
    RECT 0 866.495 0.070 866.565 ;
    RECT 0 866.635 0.070 866.705 ;
    RECT 0 866.775 0.070 866.845 ;
    RECT 0 866.915 0.070 866.985 ;
    RECT 0 867.055 0.070 867.125 ;
    RECT 0 867.195 0.070 867.265 ;
    RECT 0 867.335 0.070 867.405 ;
    RECT 0 867.475 0.070 867.545 ;
    RECT 0 867.615 0.070 867.685 ;
    RECT 0 867.755 0.070 867.825 ;
    RECT 0 867.895 0.070 867.965 ;
    RECT 0 868.035 0.070 868.105 ;
    RECT 0 868.175 0.070 868.245 ;
    RECT 0 868.315 0.070 868.385 ;
    RECT 0 868.455 0.070 868.525 ;
    RECT 0 868.595 0.070 868.665 ;
    RECT 0 868.735 0.070 868.805 ;
    RECT 0 868.875 0.070 868.945 ;
    RECT 0 869.015 0.070 869.085 ;
    RECT 0 869.155 0.070 869.225 ;
    RECT 0 869.295 0.070 869.365 ;
    RECT 0 869.435 0.070 869.505 ;
    RECT 0 869.575 0.070 869.645 ;
    RECT 0 869.715 0.070 869.785 ;
    RECT 0 869.855 0.070 869.925 ;
    RECT 0 869.995 0.070 870.065 ;
    RECT 0 870.135 0.070 870.205 ;
    RECT 0 870.275 0.070 870.345 ;
    RECT 0 870.415 0.070 870.485 ;
    RECT 0 870.555 0.070 870.625 ;
    RECT 0 870.695 0.070 870.765 ;
    RECT 0 870.835 0.070 870.905 ;
    RECT 0 870.975 0.070 871.045 ;
    RECT 0 871.115 0.070 871.185 ;
    RECT 0 871.255 0.070 871.325 ;
    RECT 0 871.395 0.070 871.465 ;
    RECT 0 871.535 0.070 871.605 ;
    RECT 0 871.675 0.070 871.745 ;
    RECT 0 871.815 0.070 871.885 ;
    RECT 0 871.955 0.070 872.025 ;
    RECT 0 872.095 0.070 872.165 ;
    RECT 0 872.235 0.070 872.305 ;
    RECT 0 872.375 0.070 872.445 ;
    RECT 0 872.515 0.070 872.585 ;
    RECT 0 872.655 0.070 872.725 ;
    RECT 0 872.795 0.070 872.865 ;
    RECT 0 872.935 0.070 873.005 ;
    RECT 0 873.075 0.070 873.145 ;
    RECT 0 873.215 0.070 873.285 ;
    RECT 0 873.355 0.070 873.425 ;
    RECT 0 873.495 0.070 873.565 ;
    RECT 0 873.635 0.070 873.705 ;
    RECT 0 873.775 0.070 873.845 ;
    RECT 0 873.915 0.070 873.985 ;
    RECT 0 874.055 0.070 874.125 ;
    RECT 0 874.195 0.070 874.265 ;
    RECT 0 874.335 0.070 874.405 ;
    RECT 0 874.475 0.070 874.545 ;
    RECT 0 874.615 0.070 874.685 ;
    RECT 0 874.755 0.070 874.825 ;
    RECT 0 874.895 0.070 874.965 ;
    RECT 0 875.035 0.070 875.105 ;
    RECT 0 875.175 0.070 875.245 ;
    RECT 0 875.315 0.070 875.385 ;
    RECT 0 875.455 0.070 875.525 ;
    RECT 0 875.595 0.070 875.665 ;
    RECT 0 875.735 0.070 875.805 ;
    RECT 0 875.875 0.070 875.945 ;
    RECT 0 876.015 0.070 876.085 ;
    RECT 0 876.155 0.070 876.225 ;
    RECT 0 876.295 0.070 876.365 ;
    RECT 0 876.435 0.070 876.505 ;
    RECT 0 876.575 0.070 876.645 ;
    RECT 0 876.715 0.070 876.785 ;
    RECT 0 876.855 0.070 876.925 ;
    RECT 0 876.995 0.070 877.065 ;
    RECT 0 877.135 0.070 877.205 ;
    RECT 0 877.275 0.070 877.345 ;
    RECT 0 877.415 0.070 877.485 ;
    RECT 0 877.555 0.070 877.625 ;
    RECT 0 877.695 0.070 877.765 ;
    RECT 0 877.835 0.070 877.905 ;
    RECT 0 877.975 0.070 878.045 ;
    RECT 0 878.115 0.070 878.185 ;
    RECT 0 878.255 0.070 878.325 ;
    RECT 0 878.395 0.070 878.465 ;
    RECT 0 878.535 0.070 878.605 ;
    RECT 0 878.675 0.070 878.745 ;
    RECT 0 878.815 0.070 878.885 ;
    RECT 0 878.955 0.070 879.025 ;
    RECT 0 879.095 0.070 879.165 ;
    RECT 0 879.235 0.070 879.305 ;
    RECT 0 879.375 0.070 879.445 ;
    RECT 0 879.515 0.070 879.585 ;
    RECT 0 879.655 0.070 879.725 ;
    RECT 0 879.795 0.070 879.865 ;
    RECT 0 879.935 0.070 880.005 ;
    RECT 0 880.075 0.070 880.145 ;
    RECT 0 880.215 0.070 880.285 ;
    RECT 0 880.355 0.070 880.425 ;
    RECT 0 880.495 0.070 880.565 ;
    RECT 0 880.635 0.070 880.705 ;
    RECT 0 880.775 0.070 880.845 ;
    RECT 0 880.915 0.070 880.985 ;
    RECT 0 881.055 0.070 881.125 ;
    RECT 0 881.195 0.070 881.265 ;
    RECT 0 881.335 0.070 881.405 ;
    RECT 0 881.475 0.070 881.545 ;
    RECT 0 881.615 0.070 881.685 ;
    RECT 0 881.755 0.070 881.825 ;
    RECT 0 881.895 0.070 881.965 ;
    RECT 0 882.035 0.070 882.105 ;
    RECT 0 882.175 0.070 882.245 ;
    RECT 0 882.315 0.070 882.385 ;
    RECT 0 882.455 0.070 882.525 ;
    RECT 0 882.595 0.070 882.665 ;
    RECT 0 882.735 0.070 882.805 ;
    RECT 0 882.875 0.070 882.945 ;
    RECT 0 883.015 0.070 883.085 ;
    RECT 0 883.155 0.070 883.225 ;
    RECT 0 883.295 0.070 883.365 ;
    RECT 0 883.435 0.070 883.505 ;
    RECT 0 883.575 0.070 883.645 ;
    RECT 0 883.715 0.070 883.785 ;
    RECT 0 883.855 0.070 883.925 ;
    RECT 0 883.995 0.070 884.065 ;
    RECT 0 884.135 0.070 884.205 ;
    RECT 0 884.275 0.070 884.345 ;
    RECT 0 884.415 0.070 884.485 ;
    RECT 0 884.555 0.070 884.625 ;
    RECT 0 884.695 0.070 884.765 ;
    RECT 0 884.835 0.070 884.905 ;
    RECT 0 884.975 0.070 885.045 ;
    RECT 0 885.115 0.070 885.185 ;
    RECT 0 885.255 0.070 885.325 ;
    RECT 0 885.395 0.070 885.465 ;
    RECT 0 885.535 0.070 885.605 ;
    RECT 0 885.675 0.070 885.745 ;
    RECT 0 885.815 0.070 885.885 ;
    RECT 0 885.955 0.070 886.025 ;
    RECT 0 886.095 0.070 886.165 ;
    RECT 0 886.235 0.070 886.305 ;
    RECT 0 886.375 0.070 886.445 ;
    RECT 0 886.515 0.070 886.585 ;
    RECT 0 886.655 0.070 886.725 ;
    RECT 0 886.795 0.070 886.865 ;
    RECT 0 886.935 0.070 887.005 ;
    RECT 0 887.075 0.070 887.145 ;
    RECT 0 887.215 0.070 887.285 ;
    RECT 0 887.355 0.070 887.425 ;
    RECT 0 887.495 0.070 887.565 ;
    RECT 0 887.635 0.070 887.705 ;
    RECT 0 887.775 0.070 887.845 ;
    RECT 0 887.915 0.070 887.985 ;
    RECT 0 888.055 0.070 888.125 ;
    RECT 0 888.195 0.070 888.265 ;
    RECT 0 888.335 0.070 888.405 ;
    RECT 0 888.475 0.070 888.545 ;
    RECT 0 888.615 0.070 888.685 ;
    RECT 0 888.755 0.070 888.825 ;
    RECT 0 888.895 0.070 888.965 ;
    RECT 0 889.035 0.070 889.105 ;
    RECT 0 889.175 0.070 889.245 ;
    RECT 0 889.315 0.070 889.385 ;
    RECT 0 889.455 0.070 889.525 ;
    RECT 0 889.595 0.070 889.665 ;
    RECT 0 889.735 0.070 889.805 ;
    RECT 0 889.875 0.070 889.945 ;
    RECT 0 890.015 0.070 890.085 ;
    RECT 0 890.155 0.070 890.225 ;
    RECT 0 890.295 0.070 890.365 ;
    RECT 0 890.435 0.070 890.505 ;
    RECT 0 890.575 0.070 890.645 ;
    RECT 0 890.715 0.070 890.785 ;
    RECT 0 890.855 0.070 890.925 ;
    RECT 0 890.995 0.070 891.065 ;
    RECT 0 891.135 0.070 891.205 ;
    RECT 0 891.275 0.070 891.345 ;
    RECT 0 891.415 0.070 891.485 ;
    RECT 0 891.555 0.070 891.625 ;
    RECT 0 891.695 0.070 891.765 ;
    RECT 0 891.835 0.070 891.905 ;
    RECT 0 891.975 0.070 892.045 ;
    RECT 0 892.115 0.070 892.185 ;
    RECT 0 892.255 0.070 892.325 ;
    RECT 0 892.395 0.070 892.465 ;
    RECT 0 892.535 0.070 892.605 ;
    RECT 0 892.675 0.070 892.745 ;
    RECT 0 892.815 0.070 892.885 ;
    RECT 0 892.955 0.070 893.025 ;
    RECT 0 893.095 0.070 893.165 ;
    RECT 0 893.235 0.070 893.305 ;
    RECT 0 893.375 0.070 893.445 ;
    RECT 0 893.515 0.070 893.585 ;
    RECT 0 893.655 0.070 893.725 ;
    RECT 0 893.795 0.070 893.865 ;
    RECT 0 893.935 0.070 894.005 ;
    RECT 0 894.075 0.070 894.145 ;
    RECT 0 894.215 0.070 894.285 ;
    RECT 0 894.355 0.070 894.425 ;
    RECT 0 894.495 0.070 894.565 ;
    RECT 0 894.635 0.070 894.705 ;
    RECT 0 894.775 0.070 894.845 ;
    RECT 0 894.915 0.070 894.985 ;
    RECT 0 895.055 0.070 895.125 ;
    RECT 0 895.195 0.070 895.265 ;
    RECT 0 895.335 0.070 895.405 ;
    RECT 0 895.475 0.070 895.545 ;
    RECT 0 895.615 0.070 895.685 ;
    RECT 0 895.755 0.070 895.825 ;
    RECT 0 895.895 0.070 895.965 ;
    RECT 0 896.035 0.070 896.105 ;
    RECT 0 896.175 0.070 896.245 ;
    RECT 0 896.315 0.070 896.385 ;
    RECT 0 896.455 0.070 896.525 ;
    RECT 0 896.595 0.070 896.665 ;
    RECT 0 896.735 0.070 896.805 ;
    RECT 0 896.875 0.070 896.945 ;
    RECT 0 897.015 0.070 897.085 ;
    RECT 0 897.155 0.070 897.225 ;
    RECT 0 897.295 0.070 897.365 ;
    RECT 0 897.435 0.070 897.505 ;
    RECT 0 897.575 0.070 897.645 ;
    RECT 0 897.715 0.070 897.785 ;
    RECT 0 897.855 0.070 897.925 ;
    RECT 0 897.995 0.070 898.065 ;
    RECT 0 898.135 0.070 898.205 ;
    RECT 0 898.275 0.070 898.345 ;
    RECT 0 898.415 0.070 898.485 ;
    RECT 0 898.555 0.070 898.625 ;
    RECT 0 898.695 0.070 898.765 ;
    RECT 0 898.835 0.070 898.905 ;
    RECT 0 898.975 0.070 899.045 ;
    RECT 0 899.115 0.070 899.185 ;
    RECT 0 899.255 0.070 899.325 ;
    RECT 0 899.395 0.070 899.465 ;
    RECT 0 899.535 0.070 899.605 ;
    RECT 0 899.675 0.070 899.745 ;
    RECT 0 899.815 0.070 899.885 ;
    RECT 0 899.955 0.070 900.025 ;
    RECT 0 900.095 0.070 900.165 ;
    RECT 0 900.235 0.070 900.305 ;
    RECT 0 900.375 0.070 900.445 ;
    RECT 0 900.515 0.070 900.585 ;
    RECT 0 900.655 0.070 900.725 ;
    RECT 0 900.795 0.070 900.865 ;
    RECT 0 900.935 0.070 901.005 ;
    RECT 0 901.075 0.070 901.145 ;
    RECT 0 901.215 0.070 901.285 ;
    RECT 0 901.355 0.070 901.425 ;
    RECT 0 901.495 0.070 901.565 ;
    RECT 0 901.635 0.070 901.705 ;
    RECT 0 901.775 0.070 901.845 ;
    RECT 0 901.915 0.070 901.985 ;
    RECT 0 902.055 0.070 902.125 ;
    RECT 0 902.195 0.070 902.265 ;
    RECT 0 902.335 0.070 902.405 ;
    RECT 0 902.475 0.070 902.545 ;
    RECT 0 902.615 0.070 902.685 ;
    RECT 0 902.755 0.070 902.825 ;
    RECT 0 902.895 0.070 902.965 ;
    RECT 0 903.035 0.070 903.105 ;
    RECT 0 903.175 0.070 1007.685 ;
    RECT 0 1007.755 0.070 1007.825 ;
    RECT 0 1007.895 0.070 1007.965 ;
    RECT 0 1008.035 0.070 1008.105 ;
    RECT 0 1008.175 0.070 1008.245 ;
    RECT 0 1008.315 0.070 1008.385 ;
    RECT 0 1008.455 0.070 1008.525 ;
    RECT 0 1008.595 0.070 1008.665 ;
    RECT 0 1008.735 0.070 1008.805 ;
    RECT 0 1008.875 0.070 1008.945 ;
    RECT 0 1009.015 0.070 1009.085 ;
    RECT 0 1009.155 0.070 1009.225 ;
    RECT 0 1009.295 0.070 1009.365 ;
    RECT 0 1009.435 0.070 1009.505 ;
    RECT 0 1009.575 0.070 1009.645 ;
    RECT 0 1009.715 0.070 1009.785 ;
    RECT 0 1009.855 0.070 1009.925 ;
    RECT 0 1009.995 0.070 1010.065 ;
    RECT 0 1010.135 0.070 1010.205 ;
    RECT 0 1010.275 0.070 1010.345 ;
    RECT 0 1010.415 0.070 1010.485 ;
    RECT 0 1010.555 0.070 1010.625 ;
    RECT 0 1010.695 0.070 1010.765 ;
    RECT 0 1010.835 0.070 1010.905 ;
    RECT 0 1010.975 0.070 1011.045 ;
    RECT 0 1011.115 0.070 1011.185 ;
    RECT 0 1011.255 0.070 1011.325 ;
    RECT 0 1011.395 0.070 1011.465 ;
    RECT 0 1011.535 0.070 1011.605 ;
    RECT 0 1011.675 0.070 1011.745 ;
    RECT 0 1011.815 0.070 1011.885 ;
    RECT 0 1011.955 0.070 1012.025 ;
    RECT 0 1012.095 0.070 1012.165 ;
    RECT 0 1012.235 0.070 1012.305 ;
    RECT 0 1012.375 0.070 1012.445 ;
    RECT 0 1012.515 0.070 1012.585 ;
    RECT 0 1012.655 0.070 1012.725 ;
    RECT 0 1012.795 0.070 1012.865 ;
    RECT 0 1012.935 0.070 1013.005 ;
    RECT 0 1013.075 0.070 1013.145 ;
    RECT 0 1013.215 0.070 1013.285 ;
    RECT 0 1013.355 0.070 1013.425 ;
    RECT 0 1013.495 0.070 1013.565 ;
    RECT 0 1013.635 0.070 1013.705 ;
    RECT 0 1013.775 0.070 1013.845 ;
    RECT 0 1013.915 0.070 1013.985 ;
    RECT 0 1014.055 0.070 1014.125 ;
    RECT 0 1014.195 0.070 1014.265 ;
    RECT 0 1014.335 0.070 1014.405 ;
    RECT 0 1014.475 0.070 1014.545 ;
    RECT 0 1014.615 0.070 1014.685 ;
    RECT 0 1014.755 0.070 1014.825 ;
    RECT 0 1014.895 0.070 1014.965 ;
    RECT 0 1015.035 0.070 1015.105 ;
    RECT 0 1015.175 0.070 1015.245 ;
    RECT 0 1015.315 0.070 1015.385 ;
    RECT 0 1015.455 0.070 1015.525 ;
    RECT 0 1015.595 0.070 1015.665 ;
    RECT 0 1015.735 0.070 1015.805 ;
    RECT 0 1015.875 0.070 1015.945 ;
    RECT 0 1016.015 0.070 1016.085 ;
    RECT 0 1016.155 0.070 1016.225 ;
    RECT 0 1016.295 0.070 1016.365 ;
    RECT 0 1016.435 0.070 1016.505 ;
    RECT 0 1016.575 0.070 1016.645 ;
    RECT 0 1016.715 0.070 1016.785 ;
    RECT 0 1016.855 0.070 1016.925 ;
    RECT 0 1016.995 0.070 1017.065 ;
    RECT 0 1017.135 0.070 1017.205 ;
    RECT 0 1017.275 0.070 1017.345 ;
    RECT 0 1017.415 0.070 1017.485 ;
    RECT 0 1017.555 0.070 1017.625 ;
    RECT 0 1017.695 0.070 1017.765 ;
    RECT 0 1017.835 0.070 1017.905 ;
    RECT 0 1017.975 0.070 1018.045 ;
    RECT 0 1018.115 0.070 1018.185 ;
    RECT 0 1018.255 0.070 1018.325 ;
    RECT 0 1018.395 0.070 1018.465 ;
    RECT 0 1018.535 0.070 1018.605 ;
    RECT 0 1018.675 0.070 1018.745 ;
    RECT 0 1018.815 0.070 1018.885 ;
    RECT 0 1018.955 0.070 1019.025 ;
    RECT 0 1019.095 0.070 1019.165 ;
    RECT 0 1019.235 0.070 1019.305 ;
    RECT 0 1019.375 0.070 1019.445 ;
    RECT 0 1019.515 0.070 1019.585 ;
    RECT 0 1019.655 0.070 1019.725 ;
    RECT 0 1019.795 0.070 1019.865 ;
    RECT 0 1019.935 0.070 1020.005 ;
    RECT 0 1020.075 0.070 1020.145 ;
    RECT 0 1020.215 0.070 1020.285 ;
    RECT 0 1020.355 0.070 1020.425 ;
    RECT 0 1020.495 0.070 1020.565 ;
    RECT 0 1020.635 0.070 1020.705 ;
    RECT 0 1020.775 0.070 1020.845 ;
    RECT 0 1020.915 0.070 1020.985 ;
    RECT 0 1021.055 0.070 1021.125 ;
    RECT 0 1021.195 0.070 1021.265 ;
    RECT 0 1021.335 0.070 1021.405 ;
    RECT 0 1021.475 0.070 1021.545 ;
    RECT 0 1021.615 0.070 1021.685 ;
    RECT 0 1021.755 0.070 1021.825 ;
    RECT 0 1021.895 0.070 1021.965 ;
    RECT 0 1022.035 0.070 1022.105 ;
    RECT 0 1022.175 0.070 1022.245 ;
    RECT 0 1022.315 0.070 1022.385 ;
    RECT 0 1022.455 0.070 1022.525 ;
    RECT 0 1022.595 0.070 1022.665 ;
    RECT 0 1022.735 0.070 1022.805 ;
    RECT 0 1022.875 0.070 1022.945 ;
    RECT 0 1023.015 0.070 1023.085 ;
    RECT 0 1023.155 0.070 1023.225 ;
    RECT 0 1023.295 0.070 1023.365 ;
    RECT 0 1023.435 0.070 1023.505 ;
    RECT 0 1023.575 0.070 1023.645 ;
    RECT 0 1023.715 0.070 1023.785 ;
    RECT 0 1023.855 0.070 1023.925 ;
    RECT 0 1023.995 0.070 1024.065 ;
    RECT 0 1024.135 0.070 1024.205 ;
    RECT 0 1024.275 0.070 1024.345 ;
    RECT 0 1024.415 0.070 1024.485 ;
    RECT 0 1024.555 0.070 1024.625 ;
    RECT 0 1024.695 0.070 1024.765 ;
    RECT 0 1024.835 0.070 1024.905 ;
    RECT 0 1024.975 0.070 1025.045 ;
    RECT 0 1025.115 0.070 1025.185 ;
    RECT 0 1025.255 0.070 1025.325 ;
    RECT 0 1025.395 0.070 1025.465 ;
    RECT 0 1025.535 0.070 1025.605 ;
    RECT 0 1025.675 0.070 1025.745 ;
    RECT 0 1025.815 0.070 1025.885 ;
    RECT 0 1025.955 0.070 1026.025 ;
    RECT 0 1026.095 0.070 1026.165 ;
    RECT 0 1026.235 0.070 1026.305 ;
    RECT 0 1026.375 0.070 1026.445 ;
    RECT 0 1026.515 0.070 1026.585 ;
    RECT 0 1026.655 0.070 1026.725 ;
    RECT 0 1026.795 0.070 1026.865 ;
    RECT 0 1026.935 0.070 1027.005 ;
    RECT 0 1027.075 0.070 1027.145 ;
    RECT 0 1027.215 0.070 1027.285 ;
    RECT 0 1027.355 0.070 1027.425 ;
    RECT 0 1027.495 0.070 1027.565 ;
    RECT 0 1027.635 0.070 1027.705 ;
    RECT 0 1027.775 0.070 1027.845 ;
    RECT 0 1027.915 0.070 1027.985 ;
    RECT 0 1028.055 0.070 1028.125 ;
    RECT 0 1028.195 0.070 1028.265 ;
    RECT 0 1028.335 0.070 1028.405 ;
    RECT 0 1028.475 0.070 1028.545 ;
    RECT 0 1028.615 0.070 1028.685 ;
    RECT 0 1028.755 0.070 1028.825 ;
    RECT 0 1028.895 0.070 1028.965 ;
    RECT 0 1029.035 0.070 1029.105 ;
    RECT 0 1029.175 0.070 1029.245 ;
    RECT 0 1029.315 0.070 1029.385 ;
    RECT 0 1029.455 0.070 1029.525 ;
    RECT 0 1029.595 0.070 1029.665 ;
    RECT 0 1029.735 0.070 1029.805 ;
    RECT 0 1029.875 0.070 1029.945 ;
    RECT 0 1030.015 0.070 1030.085 ;
    RECT 0 1030.155 0.070 1030.225 ;
    RECT 0 1030.295 0.070 1030.365 ;
    RECT 0 1030.435 0.070 1030.505 ;
    RECT 0 1030.575 0.070 1030.645 ;
    RECT 0 1030.715 0.070 1030.785 ;
    RECT 0 1030.855 0.070 1030.925 ;
    RECT 0 1030.995 0.070 1031.065 ;
    RECT 0 1031.135 0.070 1031.205 ;
    RECT 0 1031.275 0.070 1031.345 ;
    RECT 0 1031.415 0.070 1031.485 ;
    RECT 0 1031.555 0.070 1031.625 ;
    RECT 0 1031.695 0.070 1031.765 ;
    RECT 0 1031.835 0.070 1031.905 ;
    RECT 0 1031.975 0.070 1032.045 ;
    RECT 0 1032.115 0.070 1032.185 ;
    RECT 0 1032.255 0.070 1032.325 ;
    RECT 0 1032.395 0.070 1032.465 ;
    RECT 0 1032.535 0.070 1032.605 ;
    RECT 0 1032.675 0.070 1032.745 ;
    RECT 0 1032.815 0.070 1032.885 ;
    RECT 0 1032.955 0.070 1033.025 ;
    RECT 0 1033.095 0.070 1033.165 ;
    RECT 0 1033.235 0.070 1033.305 ;
    RECT 0 1033.375 0.070 1033.445 ;
    RECT 0 1033.515 0.070 1033.585 ;
    RECT 0 1033.655 0.070 1033.725 ;
    RECT 0 1033.795 0.070 1033.865 ;
    RECT 0 1033.935 0.070 1034.005 ;
    RECT 0 1034.075 0.070 1034.145 ;
    RECT 0 1034.215 0.070 1034.285 ;
    RECT 0 1034.355 0.070 1034.425 ;
    RECT 0 1034.495 0.070 1034.565 ;
    RECT 0 1034.635 0.070 1034.705 ;
    RECT 0 1034.775 0.070 1034.845 ;
    RECT 0 1034.915 0.070 1034.985 ;
    RECT 0 1035.055 0.070 1035.125 ;
    RECT 0 1035.195 0.070 1035.265 ;
    RECT 0 1035.335 0.070 1035.405 ;
    RECT 0 1035.475 0.070 1035.545 ;
    RECT 0 1035.615 0.070 1035.685 ;
    RECT 0 1035.755 0.070 1035.825 ;
    RECT 0 1035.895 0.070 1035.965 ;
    RECT 0 1036.035 0.070 1036.105 ;
    RECT 0 1036.175 0.070 1036.245 ;
    RECT 0 1036.315 0.070 1036.385 ;
    RECT 0 1036.455 0.070 1036.525 ;
    RECT 0 1036.595 0.070 1036.665 ;
    RECT 0 1036.735 0.070 1036.805 ;
    RECT 0 1036.875 0.070 1036.945 ;
    RECT 0 1037.015 0.070 1037.085 ;
    RECT 0 1037.155 0.070 1037.225 ;
    RECT 0 1037.295 0.070 1037.365 ;
    RECT 0 1037.435 0.070 1037.505 ;
    RECT 0 1037.575 0.070 1037.645 ;
    RECT 0 1037.715 0.070 1037.785 ;
    RECT 0 1037.855 0.070 1037.925 ;
    RECT 0 1037.995 0.070 1038.065 ;
    RECT 0 1038.135 0.070 1038.205 ;
    RECT 0 1038.275 0.070 1038.345 ;
    RECT 0 1038.415 0.070 1038.485 ;
    RECT 0 1038.555 0.070 1038.625 ;
    RECT 0 1038.695 0.070 1038.765 ;
    RECT 0 1038.835 0.070 1038.905 ;
    RECT 0 1038.975 0.070 1039.045 ;
    RECT 0 1039.115 0.070 1039.185 ;
    RECT 0 1039.255 0.070 1039.325 ;
    RECT 0 1039.395 0.070 1039.465 ;
    RECT 0 1039.535 0.070 1039.605 ;
    RECT 0 1039.675 0.070 1039.745 ;
    RECT 0 1039.815 0.070 1039.885 ;
    RECT 0 1039.955 0.070 1040.025 ;
    RECT 0 1040.095 0.070 1040.165 ;
    RECT 0 1040.235 0.070 1040.305 ;
    RECT 0 1040.375 0.070 1040.445 ;
    RECT 0 1040.515 0.070 1040.585 ;
    RECT 0 1040.655 0.070 1040.725 ;
    RECT 0 1040.795 0.070 1040.865 ;
    RECT 0 1040.935 0.070 1041.005 ;
    RECT 0 1041.075 0.070 1041.145 ;
    RECT 0 1041.215 0.070 1041.285 ;
    RECT 0 1041.355 0.070 1041.425 ;
    RECT 0 1041.495 0.070 1041.565 ;
    RECT 0 1041.635 0.070 1041.705 ;
    RECT 0 1041.775 0.070 1041.845 ;
    RECT 0 1041.915 0.070 1041.985 ;
    RECT 0 1042.055 0.070 1042.125 ;
    RECT 0 1042.195 0.070 1042.265 ;
    RECT 0 1042.335 0.070 1042.405 ;
    RECT 0 1042.475 0.070 1042.545 ;
    RECT 0 1042.615 0.070 1042.685 ;
    RECT 0 1042.755 0.070 1042.825 ;
    RECT 0 1042.895 0.070 1042.965 ;
    RECT 0 1043.035 0.070 1043.105 ;
    RECT 0 1043.175 0.070 1043.245 ;
    RECT 0 1043.315 0.070 1043.385 ;
    RECT 0 1043.455 0.070 1043.525 ;
    RECT 0 1043.595 0.070 1043.665 ;
    RECT 0 1043.735 0.070 1043.805 ;
    RECT 0 1043.875 0.070 1043.945 ;
    RECT 0 1044.015 0.070 1044.085 ;
    RECT 0 1044.155 0.070 1044.225 ;
    RECT 0 1044.295 0.070 1044.365 ;
    RECT 0 1044.435 0.070 1044.505 ;
    RECT 0 1044.575 0.070 1044.645 ;
    RECT 0 1044.715 0.070 1044.785 ;
    RECT 0 1044.855 0.070 1044.925 ;
    RECT 0 1044.995 0.070 1045.065 ;
    RECT 0 1045.135 0.070 1045.205 ;
    RECT 0 1045.275 0.070 1045.345 ;
    RECT 0 1045.415 0.070 1045.485 ;
    RECT 0 1045.555 0.070 1045.625 ;
    RECT 0 1045.695 0.070 1045.765 ;
    RECT 0 1045.835 0.070 1045.905 ;
    RECT 0 1045.975 0.070 1046.045 ;
    RECT 0 1046.115 0.070 1046.185 ;
    RECT 0 1046.255 0.070 1046.325 ;
    RECT 0 1046.395 0.070 1046.465 ;
    RECT 0 1046.535 0.070 1046.605 ;
    RECT 0 1046.675 0.070 1046.745 ;
    RECT 0 1046.815 0.070 1046.885 ;
    RECT 0 1046.955 0.070 1047.025 ;
    RECT 0 1047.095 0.070 1047.165 ;
    RECT 0 1047.235 0.070 1047.305 ;
    RECT 0 1047.375 0.070 1047.445 ;
    RECT 0 1047.515 0.070 1047.585 ;
    RECT 0 1047.655 0.070 1047.725 ;
    RECT 0 1047.795 0.070 1047.865 ;
    RECT 0 1047.935 0.070 1048.005 ;
    RECT 0 1048.075 0.070 1048.145 ;
    RECT 0 1048.215 0.070 1048.285 ;
    RECT 0 1048.355 0.070 1048.425 ;
    RECT 0 1048.495 0.070 1048.565 ;
    RECT 0 1048.635 0.070 1048.705 ;
    RECT 0 1048.775 0.070 1048.845 ;
    RECT 0 1048.915 0.070 1048.985 ;
    RECT 0 1049.055 0.070 1049.125 ;
    RECT 0 1049.195 0.070 1049.265 ;
    RECT 0 1049.335 0.070 1049.405 ;
    RECT 0 1049.475 0.070 1049.545 ;
    RECT 0 1049.615 0.070 1049.685 ;
    RECT 0 1049.755 0.070 1049.825 ;
    RECT 0 1049.895 0.070 1049.965 ;
    RECT 0 1050.035 0.070 1050.105 ;
    RECT 0 1050.175 0.070 1050.245 ;
    RECT 0 1050.315 0.070 1050.385 ;
    RECT 0 1050.455 0.070 1050.525 ;
    RECT 0 1050.595 0.070 1050.665 ;
    RECT 0 1050.735 0.070 1050.805 ;
    RECT 0 1050.875 0.070 1050.945 ;
    RECT 0 1051.015 0.070 1051.085 ;
    RECT 0 1051.155 0.070 1051.225 ;
    RECT 0 1051.295 0.070 1051.365 ;
    RECT 0 1051.435 0.070 1051.505 ;
    RECT 0 1051.575 0.070 1051.645 ;
    RECT 0 1051.715 0.070 1051.785 ;
    RECT 0 1051.855 0.070 1051.925 ;
    RECT 0 1051.995 0.070 1052.065 ;
    RECT 0 1052.135 0.070 1052.205 ;
    RECT 0 1052.275 0.070 1052.345 ;
    RECT 0 1052.415 0.070 1052.485 ;
    RECT 0 1052.555 0.070 1052.625 ;
    RECT 0 1052.695 0.070 1052.765 ;
    RECT 0 1052.835 0.070 1052.905 ;
    RECT 0 1052.975 0.070 1053.045 ;
    RECT 0 1053.115 0.070 1053.185 ;
    RECT 0 1053.255 0.070 1053.325 ;
    RECT 0 1053.395 0.070 1053.465 ;
    RECT 0 1053.535 0.070 1053.605 ;
    RECT 0 1053.675 0.070 1053.745 ;
    RECT 0 1053.815 0.070 1053.885 ;
    RECT 0 1053.955 0.070 1054.025 ;
    RECT 0 1054.095 0.070 1054.165 ;
    RECT 0 1054.235 0.070 1054.305 ;
    RECT 0 1054.375 0.070 1054.445 ;
    RECT 0 1054.515 0.070 1054.585 ;
    RECT 0 1054.655 0.070 1054.725 ;
    RECT 0 1054.795 0.070 1054.865 ;
    RECT 0 1054.935 0.070 1055.005 ;
    RECT 0 1055.075 0.070 1055.145 ;
    RECT 0 1055.215 0.070 1055.285 ;
    RECT 0 1055.355 0.070 1055.425 ;
    RECT 0 1055.495 0.070 1055.565 ;
    RECT 0 1055.635 0.070 1055.705 ;
    RECT 0 1055.775 0.070 1055.845 ;
    RECT 0 1055.915 0.070 1055.985 ;
    RECT 0 1056.055 0.070 1056.125 ;
    RECT 0 1056.195 0.070 1056.265 ;
    RECT 0 1056.335 0.070 1056.405 ;
    RECT 0 1056.475 0.070 1056.545 ;
    RECT 0 1056.615 0.070 1056.685 ;
    RECT 0 1056.755 0.070 1056.825 ;
    RECT 0 1056.895 0.070 1056.965 ;
    RECT 0 1057.035 0.070 1057.105 ;
    RECT 0 1057.175 0.070 1057.245 ;
    RECT 0 1057.315 0.070 1057.385 ;
    RECT 0 1057.455 0.070 1057.525 ;
    RECT 0 1057.595 0.070 1057.665 ;
    RECT 0 1057.735 0.070 1057.805 ;
    RECT 0 1057.875 0.070 1057.945 ;
    RECT 0 1058.015 0.070 1058.085 ;
    RECT 0 1058.155 0.070 1058.225 ;
    RECT 0 1058.295 0.070 1058.365 ;
    RECT 0 1058.435 0.070 1058.505 ;
    RECT 0 1058.575 0.070 1058.645 ;
    RECT 0 1058.715 0.070 1058.785 ;
    RECT 0 1058.855 0.070 1058.925 ;
    RECT 0 1058.995 0.070 1059.065 ;
    RECT 0 1059.135 0.070 1059.205 ;
    RECT 0 1059.275 0.070 1059.345 ;
    RECT 0 1059.415 0.070 1059.485 ;
    RECT 0 1059.555 0.070 1059.625 ;
    RECT 0 1059.695 0.070 1059.765 ;
    RECT 0 1059.835 0.070 1059.905 ;
    RECT 0 1059.975 0.070 1060.045 ;
    RECT 0 1060.115 0.070 1060.185 ;
    RECT 0 1060.255 0.070 1060.325 ;
    RECT 0 1060.395 0.070 1060.465 ;
    RECT 0 1060.535 0.070 1060.605 ;
    RECT 0 1060.675 0.070 1060.745 ;
    RECT 0 1060.815 0.070 1060.885 ;
    RECT 0 1060.955 0.070 1061.025 ;
    RECT 0 1061.095 0.070 1061.165 ;
    RECT 0 1061.235 0.070 1061.305 ;
    RECT 0 1061.375 0.070 1061.445 ;
    RECT 0 1061.515 0.070 1061.585 ;
    RECT 0 1061.655 0.070 1061.725 ;
    RECT 0 1061.795 0.070 1061.865 ;
    RECT 0 1061.935 0.070 1062.005 ;
    RECT 0 1062.075 0.070 1062.145 ;
    RECT 0 1062.215 0.070 1062.285 ;
    RECT 0 1062.355 0.070 1062.425 ;
    RECT 0 1062.495 0.070 1062.565 ;
    RECT 0 1062.635 0.070 1062.705 ;
    RECT 0 1062.775 0.070 1062.845 ;
    RECT 0 1062.915 0.070 1062.985 ;
    RECT 0 1063.055 0.070 1063.125 ;
    RECT 0 1063.195 0.070 1063.265 ;
    RECT 0 1063.335 0.070 1063.405 ;
    RECT 0 1063.475 0.070 1063.545 ;
    RECT 0 1063.615 0.070 1063.685 ;
    RECT 0 1063.755 0.070 1063.825 ;
    RECT 0 1063.895 0.070 1063.965 ;
    RECT 0 1064.035 0.070 1064.105 ;
    RECT 0 1064.175 0.070 1064.245 ;
    RECT 0 1064.315 0.070 1064.385 ;
    RECT 0 1064.455 0.070 1064.525 ;
    RECT 0 1064.595 0.070 1064.665 ;
    RECT 0 1064.735 0.070 1064.805 ;
    RECT 0 1064.875 0.070 1064.945 ;
    RECT 0 1065.015 0.070 1065.085 ;
    RECT 0 1065.155 0.070 1065.225 ;
    RECT 0 1065.295 0.070 1065.365 ;
    RECT 0 1065.435 0.070 1065.505 ;
    RECT 0 1065.575 0.070 1065.645 ;
    RECT 0 1065.715 0.070 1065.785 ;
    RECT 0 1065.855 0.070 1065.925 ;
    RECT 0 1065.995 0.070 1066.065 ;
    RECT 0 1066.135 0.070 1066.205 ;
    RECT 0 1066.275 0.070 1066.345 ;
    RECT 0 1066.415 0.070 1066.485 ;
    RECT 0 1066.555 0.070 1066.625 ;
    RECT 0 1066.695 0.070 1066.765 ;
    RECT 0 1066.835 0.070 1066.905 ;
    RECT 0 1066.975 0.070 1067.045 ;
    RECT 0 1067.115 0.070 1067.185 ;
    RECT 0 1067.255 0.070 1067.325 ;
    RECT 0 1067.395 0.070 1067.465 ;
    RECT 0 1067.535 0.070 1067.605 ;
    RECT 0 1067.675 0.070 1067.745 ;
    RECT 0 1067.815 0.070 1067.885 ;
    RECT 0 1067.955 0.070 1068.025 ;
    RECT 0 1068.095 0.070 1068.165 ;
    RECT 0 1068.235 0.070 1068.305 ;
    RECT 0 1068.375 0.070 1068.445 ;
    RECT 0 1068.515 0.070 1068.585 ;
    RECT 0 1068.655 0.070 1068.725 ;
    RECT 0 1068.795 0.070 1068.865 ;
    RECT 0 1068.935 0.070 1069.005 ;
    RECT 0 1069.075 0.070 1069.145 ;
    RECT 0 1069.215 0.070 1069.285 ;
    RECT 0 1069.355 0.070 1069.425 ;
    RECT 0 1069.495 0.070 1069.565 ;
    RECT 0 1069.635 0.070 1069.705 ;
    RECT 0 1069.775 0.070 1069.845 ;
    RECT 0 1069.915 0.070 1069.985 ;
    RECT 0 1070.055 0.070 1070.125 ;
    RECT 0 1070.195 0.070 1070.265 ;
    RECT 0 1070.335 0.070 1070.405 ;
    RECT 0 1070.475 0.070 1070.545 ;
    RECT 0 1070.615 0.070 1070.685 ;
    RECT 0 1070.755 0.070 1070.825 ;
    RECT 0 1070.895 0.070 1070.965 ;
    RECT 0 1071.035 0.070 1071.105 ;
    RECT 0 1071.175 0.070 1071.245 ;
    RECT 0 1071.315 0.070 1071.385 ;
    RECT 0 1071.455 0.070 1071.525 ;
    RECT 0 1071.595 0.070 1071.665 ;
    RECT 0 1071.735 0.070 1071.805 ;
    RECT 0 1071.875 0.070 1071.945 ;
    RECT 0 1072.015 0.070 1072.085 ;
    RECT 0 1072.155 0.070 1072.225 ;
    RECT 0 1072.295 0.070 1072.365 ;
    RECT 0 1072.435 0.070 1072.505 ;
    RECT 0 1072.575 0.070 1072.645 ;
    RECT 0 1072.715 0.070 1072.785 ;
    RECT 0 1072.855 0.070 1072.925 ;
    RECT 0 1072.995 0.070 1073.065 ;
    RECT 0 1073.135 0.070 1073.205 ;
    RECT 0 1073.275 0.070 1073.345 ;
    RECT 0 1073.415 0.070 1073.485 ;
    RECT 0 1073.555 0.070 1073.625 ;
    RECT 0 1073.695 0.070 1073.765 ;
    RECT 0 1073.835 0.070 1073.905 ;
    RECT 0 1073.975 0.070 1074.045 ;
    RECT 0 1074.115 0.070 1074.185 ;
    RECT 0 1074.255 0.070 1074.325 ;
    RECT 0 1074.395 0.070 1074.465 ;
    RECT 0 1074.535 0.070 1074.605 ;
    RECT 0 1074.675 0.070 1074.745 ;
    RECT 0 1074.815 0.070 1074.885 ;
    RECT 0 1074.955 0.070 1075.025 ;
    RECT 0 1075.095 0.070 1075.165 ;
    RECT 0 1075.235 0.070 1075.305 ;
    RECT 0 1075.375 0.070 1075.445 ;
    RECT 0 1075.515 0.070 1075.585 ;
    RECT 0 1075.655 0.070 1075.725 ;
    RECT 0 1075.795 0.070 1075.865 ;
    RECT 0 1075.935 0.070 1076.005 ;
    RECT 0 1076.075 0.070 1076.145 ;
    RECT 0 1076.215 0.070 1076.285 ;
    RECT 0 1076.355 0.070 1076.425 ;
    RECT 0 1076.495 0.070 1076.565 ;
    RECT 0 1076.635 0.070 1076.705 ;
    RECT 0 1076.775 0.070 1076.845 ;
    RECT 0 1076.915 0.070 1076.985 ;
    RECT 0 1077.055 0.070 1077.125 ;
    RECT 0 1077.195 0.070 1077.265 ;
    RECT 0 1077.335 0.070 1077.405 ;
    RECT 0 1077.475 0.070 1077.545 ;
    RECT 0 1077.615 0.070 1077.685 ;
    RECT 0 1077.755 0.070 1077.825 ;
    RECT 0 1077.895 0.070 1077.965 ;
    RECT 0 1078.035 0.070 1078.105 ;
    RECT 0 1078.175 0.070 1078.245 ;
    RECT 0 1078.315 0.070 1078.385 ;
    RECT 0 1078.455 0.070 1078.525 ;
    RECT 0 1078.595 0.070 1078.665 ;
    RECT 0 1078.735 0.070 1078.805 ;
    RECT 0 1078.875 0.070 1078.945 ;
    RECT 0 1079.015 0.070 1079.085 ;
    RECT 0 1079.155 0.070 1079.225 ;
    RECT 0 1079.295 0.070 1079.365 ;
    RECT 0 1079.435 0.070 1079.505 ;
    RECT 0 1079.575 0.070 1079.645 ;
    RECT 0 1079.715 0.070 1079.785 ;
    RECT 0 1079.855 0.070 1079.925 ;
    RECT 0 1079.995 0.070 1080.065 ;
    RECT 0 1080.135 0.070 1080.205 ;
    RECT 0 1080.275 0.070 1080.345 ;
    RECT 0 1080.415 0.070 1080.485 ;
    RECT 0 1080.555 0.070 1080.625 ;
    RECT 0 1080.695 0.070 1080.765 ;
    RECT 0 1080.835 0.070 1080.905 ;
    RECT 0 1080.975 0.070 1081.045 ;
    RECT 0 1081.115 0.070 1081.185 ;
    RECT 0 1081.255 0.070 1081.325 ;
    RECT 0 1081.395 0.070 1081.465 ;
    RECT 0 1081.535 0.070 1081.605 ;
    RECT 0 1081.675 0.070 1081.745 ;
    RECT 0 1081.815 0.070 1081.885 ;
    RECT 0 1081.955 0.070 1082.025 ;
    RECT 0 1082.095 0.070 1082.165 ;
    RECT 0 1082.235 0.070 1082.305 ;
    RECT 0 1082.375 0.070 1082.445 ;
    RECT 0 1082.515 0.070 1082.585 ;
    RECT 0 1082.655 0.070 1082.725 ;
    RECT 0 1082.795 0.070 1082.865 ;
    RECT 0 1082.935 0.070 1083.005 ;
    RECT 0 1083.075 0.070 1083.145 ;
    RECT 0 1083.215 0.070 1083.285 ;
    RECT 0 1083.355 0.070 1083.425 ;
    RECT 0 1083.495 0.070 1083.565 ;
    RECT 0 1083.635 0.070 1083.705 ;
    RECT 0 1083.775 0.070 1083.845 ;
    RECT 0 1083.915 0.070 1083.985 ;
    RECT 0 1084.055 0.070 1084.125 ;
    RECT 0 1084.195 0.070 1084.265 ;
    RECT 0 1084.335 0.070 1084.405 ;
    RECT 0 1084.475 0.070 1084.545 ;
    RECT 0 1084.615 0.070 1084.685 ;
    RECT 0 1084.755 0.070 1084.825 ;
    RECT 0 1084.895 0.070 1084.965 ;
    RECT 0 1085.035 0.070 1085.105 ;
    RECT 0 1085.175 0.070 1085.245 ;
    RECT 0 1085.315 0.070 1085.385 ;
    RECT 0 1085.455 0.070 1085.525 ;
    RECT 0 1085.595 0.070 1085.665 ;
    RECT 0 1085.735 0.070 1085.805 ;
    RECT 0 1085.875 0.070 1085.945 ;
    RECT 0 1086.015 0.070 1086.085 ;
    RECT 0 1086.155 0.070 1086.225 ;
    RECT 0 1086.295 0.070 1086.365 ;
    RECT 0 1086.435 0.070 1086.505 ;
    RECT 0 1086.575 0.070 1086.645 ;
    RECT 0 1086.715 0.070 1086.785 ;
    RECT 0 1086.855 0.070 1086.925 ;
    RECT 0 1086.995 0.070 1087.065 ;
    RECT 0 1087.135 0.070 1087.205 ;
    RECT 0 1087.275 0.070 1087.345 ;
    RECT 0 1087.415 0.070 1087.485 ;
    RECT 0 1087.555 0.070 1087.625 ;
    RECT 0 1087.695 0.070 1087.765 ;
    RECT 0 1087.835 0.070 1087.905 ;
    RECT 0 1087.975 0.070 1088.045 ;
    RECT 0 1088.115 0.070 1088.185 ;
    RECT 0 1088.255 0.070 1088.325 ;
    RECT 0 1088.395 0.070 1088.465 ;
    RECT 0 1088.535 0.070 1088.605 ;
    RECT 0 1088.675 0.070 1088.745 ;
    RECT 0 1088.815 0.070 1088.885 ;
    RECT 0 1088.955 0.070 1089.025 ;
    RECT 0 1089.095 0.070 1089.165 ;
    RECT 0 1089.235 0.070 1089.305 ;
    RECT 0 1089.375 0.070 1089.445 ;
    RECT 0 1089.515 0.070 1089.585 ;
    RECT 0 1089.655 0.070 1089.725 ;
    RECT 0 1089.795 0.070 1089.865 ;
    RECT 0 1089.935 0.070 1090.005 ;
    RECT 0 1090.075 0.070 1090.145 ;
    RECT 0 1090.215 0.070 1090.285 ;
    RECT 0 1090.355 0.070 1090.425 ;
    RECT 0 1090.495 0.070 1090.565 ;
    RECT 0 1090.635 0.070 1090.705 ;
    RECT 0 1090.775 0.070 1090.845 ;
    RECT 0 1090.915 0.070 1090.985 ;
    RECT 0 1091.055 0.070 1091.125 ;
    RECT 0 1091.195 0.070 1091.265 ;
    RECT 0 1091.335 0.070 1091.405 ;
    RECT 0 1091.475 0.070 1091.545 ;
    RECT 0 1091.615 0.070 1091.685 ;
    RECT 0 1091.755 0.070 1091.825 ;
    RECT 0 1091.895 0.070 1091.965 ;
    RECT 0 1092.035 0.070 1092.105 ;
    RECT 0 1092.175 0.070 1092.245 ;
    RECT 0 1092.315 0.070 1092.385 ;
    RECT 0 1092.455 0.070 1092.525 ;
    RECT 0 1092.595 0.070 1092.665 ;
    RECT 0 1092.735 0.070 1092.805 ;
    RECT 0 1092.875 0.070 1092.945 ;
    RECT 0 1093.015 0.070 1093.085 ;
    RECT 0 1093.155 0.070 1093.225 ;
    RECT 0 1093.295 0.070 1093.365 ;
    RECT 0 1093.435 0.070 1093.505 ;
    RECT 0 1093.575 0.070 1093.645 ;
    RECT 0 1093.715 0.070 1093.785 ;
    RECT 0 1093.855 0.070 1093.925 ;
    RECT 0 1093.995 0.070 1094.065 ;
    RECT 0 1094.135 0.070 1094.205 ;
    RECT 0 1094.275 0.070 1094.345 ;
    RECT 0 1094.415 0.070 1094.485 ;
    RECT 0 1094.555 0.070 1094.625 ;
    RECT 0 1094.695 0.070 1094.765 ;
    RECT 0 1094.835 0.070 1094.905 ;
    RECT 0 1094.975 0.070 1095.045 ;
    RECT 0 1095.115 0.070 1095.185 ;
    RECT 0 1095.255 0.070 1095.325 ;
    RECT 0 1095.395 0.070 1095.465 ;
    RECT 0 1095.535 0.070 1095.605 ;
    RECT 0 1095.675 0.070 1095.745 ;
    RECT 0 1095.815 0.070 1095.885 ;
    RECT 0 1095.955 0.070 1096.025 ;
    RECT 0 1096.095 0.070 1096.165 ;
    RECT 0 1096.235 0.070 1096.305 ;
    RECT 0 1096.375 0.070 1096.445 ;
    RECT 0 1096.515 0.070 1096.585 ;
    RECT 0 1096.655 0.070 1096.725 ;
    RECT 0 1096.795 0.070 1096.865 ;
    RECT 0 1096.935 0.070 1097.005 ;
    RECT 0 1097.075 0.070 1097.145 ;
    RECT 0 1097.215 0.070 1097.285 ;
    RECT 0 1097.355 0.070 1097.425 ;
    RECT 0 1097.495 0.070 1097.565 ;
    RECT 0 1097.635 0.070 1097.705 ;
    RECT 0 1097.775 0.070 1097.845 ;
    RECT 0 1097.915 0.070 1097.985 ;
    RECT 0 1098.055 0.070 1098.125 ;
    RECT 0 1098.195 0.070 1098.265 ;
    RECT 0 1098.335 0.070 1098.405 ;
    RECT 0 1098.475 0.070 1098.545 ;
    RECT 0 1098.615 0.070 1098.685 ;
    RECT 0 1098.755 0.070 1098.825 ;
    RECT 0 1098.895 0.070 1098.965 ;
    RECT 0 1099.035 0.070 1099.105 ;
    RECT 0 1099.175 0.070 1099.245 ;
    RECT 0 1099.315 0.070 1099.385 ;
    RECT 0 1099.455 0.070 1099.525 ;
    RECT 0 1099.595 0.070 1099.665 ;
    RECT 0 1099.735 0.070 1099.805 ;
    RECT 0 1099.875 0.070 1099.945 ;
    RECT 0 1100.015 0.070 1100.085 ;
    RECT 0 1100.155 0.070 1100.225 ;
    RECT 0 1100.295 0.070 1100.365 ;
    RECT 0 1100.435 0.070 1100.505 ;
    RECT 0 1100.575 0.070 1100.645 ;
    RECT 0 1100.715 0.070 1100.785 ;
    RECT 0 1100.855 0.070 1100.925 ;
    RECT 0 1100.995 0.070 1101.065 ;
    RECT 0 1101.135 0.070 1101.205 ;
    RECT 0 1101.275 0.070 1101.345 ;
    RECT 0 1101.415 0.070 1101.485 ;
    RECT 0 1101.555 0.070 1101.625 ;
    RECT 0 1101.695 0.070 1101.765 ;
    RECT 0 1101.835 0.070 1101.905 ;
    RECT 0 1101.975 0.070 1102.045 ;
    RECT 0 1102.115 0.070 1102.185 ;
    RECT 0 1102.255 0.070 1102.325 ;
    RECT 0 1102.395 0.070 1102.465 ;
    RECT 0 1102.535 0.070 1102.605 ;
    RECT 0 1102.675 0.070 1102.745 ;
    RECT 0 1102.815 0.070 1102.885 ;
    RECT 0 1102.955 0.070 1103.025 ;
    RECT 0 1103.095 0.070 1103.165 ;
    RECT 0 1103.235 0.070 1103.305 ;
    RECT 0 1103.375 0.070 1103.445 ;
    RECT 0 1103.515 0.070 1103.585 ;
    RECT 0 1103.655 0.070 1103.725 ;
    RECT 0 1103.795 0.070 1103.865 ;
    RECT 0 1103.935 0.070 1104.005 ;
    RECT 0 1104.075 0.070 1104.145 ;
    RECT 0 1104.215 0.070 1104.285 ;
    RECT 0 1104.355 0.070 1104.425 ;
    RECT 0 1104.495 0.070 1104.565 ;
    RECT 0 1104.635 0.070 1104.705 ;
    RECT 0 1104.775 0.070 1104.845 ;
    RECT 0 1104.915 0.070 1104.985 ;
    RECT 0 1105.055 0.070 1105.125 ;
    RECT 0 1105.195 0.070 1105.265 ;
    RECT 0 1105.335 0.070 1105.405 ;
    RECT 0 1105.475 0.070 1105.545 ;
    RECT 0 1105.615 0.070 1105.685 ;
    RECT 0 1105.755 0.070 1105.825 ;
    RECT 0 1105.895 0.070 1105.965 ;
    RECT 0 1106.035 0.070 1106.105 ;
    RECT 0 1106.175 0.070 1106.245 ;
    RECT 0 1106.315 0.070 1106.385 ;
    RECT 0 1106.455 0.070 1106.525 ;
    RECT 0 1106.595 0.070 1106.665 ;
    RECT 0 1106.735 0.070 1106.805 ;
    RECT 0 1106.875 0.070 1106.945 ;
    RECT 0 1107.015 0.070 1107.085 ;
    RECT 0 1107.155 0.070 1107.225 ;
    RECT 0 1107.295 0.070 1107.365 ;
    RECT 0 1107.435 0.070 1107.505 ;
    RECT 0 1107.575 0.070 1107.645 ;
    RECT 0 1107.715 0.070 1107.785 ;
    RECT 0 1107.855 0.070 1107.925 ;
    RECT 0 1107.995 0.070 1108.065 ;
    RECT 0 1108.135 0.070 1108.205 ;
    RECT 0 1108.275 0.070 1108.345 ;
    RECT 0 1108.415 0.070 1108.485 ;
    RECT 0 1108.555 0.070 1108.625 ;
    RECT 0 1108.695 0.070 1108.765 ;
    RECT 0 1108.835 0.070 1108.905 ;
    RECT 0 1108.975 0.070 1109.045 ;
    RECT 0 1109.115 0.070 1109.185 ;
    RECT 0 1109.255 0.070 1109.325 ;
    RECT 0 1109.395 0.070 1109.465 ;
    RECT 0 1109.535 0.070 1109.605 ;
    RECT 0 1109.675 0.070 1109.745 ;
    RECT 0 1109.815 0.070 1109.885 ;
    RECT 0 1109.955 0.070 1110.025 ;
    RECT 0 1110.095 0.070 1110.165 ;
    RECT 0 1110.235 0.070 1110.305 ;
    RECT 0 1110.375 0.070 1110.445 ;
    RECT 0 1110.515 0.070 1110.585 ;
    RECT 0 1110.655 0.070 1110.725 ;
    RECT 0 1110.795 0.070 1110.865 ;
    RECT 0 1110.935 0.070 1111.005 ;
    RECT 0 1111.075 0.070 1111.145 ;
    RECT 0 1111.215 0.070 1111.285 ;
    RECT 0 1111.355 0.070 1111.425 ;
    RECT 0 1111.495 0.070 1111.565 ;
    RECT 0 1111.635 0.070 1111.705 ;
    RECT 0 1111.775 0.070 1111.845 ;
    RECT 0 1111.915 0.070 1111.985 ;
    RECT 0 1112.055 0.070 1112.125 ;
    RECT 0 1112.195 0.070 1112.265 ;
    RECT 0 1112.335 0.070 1112.405 ;
    RECT 0 1112.475 0.070 1112.545 ;
    RECT 0 1112.615 0.070 1112.685 ;
    RECT 0 1112.755 0.070 1112.825 ;
    RECT 0 1112.895 0.070 1112.965 ;
    RECT 0 1113.035 0.070 1113.105 ;
    RECT 0 1113.175 0.070 1113.245 ;
    RECT 0 1113.315 0.070 1113.385 ;
    RECT 0 1113.455 0.070 1113.525 ;
    RECT 0 1113.595 0.070 1113.665 ;
    RECT 0 1113.735 0.070 1113.805 ;
    RECT 0 1113.875 0.070 1113.945 ;
    RECT 0 1114.015 0.070 1114.085 ;
    RECT 0 1114.155 0.070 1114.225 ;
    RECT 0 1114.295 0.070 1114.365 ;
    RECT 0 1114.435 0.070 1114.505 ;
    RECT 0 1114.575 0.070 1114.645 ;
    RECT 0 1114.715 0.070 1114.785 ;
    RECT 0 1114.855 0.070 1114.925 ;
    RECT 0 1114.995 0.070 1115.065 ;
    RECT 0 1115.135 0.070 1115.205 ;
    RECT 0 1115.275 0.070 1115.345 ;
    RECT 0 1115.415 0.070 1115.485 ;
    RECT 0 1115.555 0.070 1115.625 ;
    RECT 0 1115.695 0.070 1115.765 ;
    RECT 0 1115.835 0.070 1115.905 ;
    RECT 0 1115.975 0.070 1116.045 ;
    RECT 0 1116.115 0.070 1116.185 ;
    RECT 0 1116.255 0.070 1116.325 ;
    RECT 0 1116.395 0.070 1116.465 ;
    RECT 0 1116.535 0.070 1116.605 ;
    RECT 0 1116.675 0.070 1116.745 ;
    RECT 0 1116.815 0.070 1116.885 ;
    RECT 0 1116.955 0.070 1117.025 ;
    RECT 0 1117.095 0.070 1117.165 ;
    RECT 0 1117.235 0.070 1117.305 ;
    RECT 0 1117.375 0.070 1117.445 ;
    RECT 0 1117.515 0.070 1117.585 ;
    RECT 0 1117.655 0.070 1117.725 ;
    RECT 0 1117.795 0.070 1117.865 ;
    RECT 0 1117.935 0.070 1118.005 ;
    RECT 0 1118.075 0.070 1118.145 ;
    RECT 0 1118.215 0.070 1118.285 ;
    RECT 0 1118.355 0.070 1118.425 ;
    RECT 0 1118.495 0.070 1118.565 ;
    RECT 0 1118.635 0.070 1118.705 ;
    RECT 0 1118.775 0.070 1118.845 ;
    RECT 0 1118.915 0.070 1118.985 ;
    RECT 0 1119.055 0.070 1119.125 ;
    RECT 0 1119.195 0.070 1119.265 ;
    RECT 0 1119.335 0.070 1119.405 ;
    RECT 0 1119.475 0.070 1119.545 ;
    RECT 0 1119.615 0.070 1119.685 ;
    RECT 0 1119.755 0.070 1119.825 ;
    RECT 0 1119.895 0.070 1119.965 ;
    RECT 0 1120.035 0.070 1120.105 ;
    RECT 0 1120.175 0.070 1120.245 ;
    RECT 0 1120.315 0.070 1120.385 ;
    RECT 0 1120.455 0.070 1120.525 ;
    RECT 0 1120.595 0.070 1120.665 ;
    RECT 0 1120.735 0.070 1120.805 ;
    RECT 0 1120.875 0.070 1120.945 ;
    RECT 0 1121.015 0.070 1121.085 ;
    RECT 0 1121.155 0.070 1121.225 ;
    RECT 0 1121.295 0.070 1121.365 ;
    RECT 0 1121.435 0.070 1121.505 ;
    RECT 0 1121.575 0.070 1121.645 ;
    RECT 0 1121.715 0.070 1121.785 ;
    RECT 0 1121.855 0.070 1121.925 ;
    RECT 0 1121.995 0.070 1122.065 ;
    RECT 0 1122.135 0.070 1122.205 ;
    RECT 0 1122.275 0.070 1122.345 ;
    RECT 0 1122.415 0.070 1122.485 ;
    RECT 0 1122.555 0.070 1122.625 ;
    RECT 0 1122.695 0.070 1122.765 ;
    RECT 0 1122.835 0.070 1122.905 ;
    RECT 0 1122.975 0.070 1123.045 ;
    RECT 0 1123.115 0.070 1123.185 ;
    RECT 0 1123.255 0.070 1123.325 ;
    RECT 0 1123.395 0.070 1123.465 ;
    RECT 0 1123.535 0.070 1123.605 ;
    RECT 0 1123.675 0.070 1123.745 ;
    RECT 0 1123.815 0.070 1123.885 ;
    RECT 0 1123.955 0.070 1124.025 ;
    RECT 0 1124.095 0.070 1124.165 ;
    RECT 0 1124.235 0.070 1124.305 ;
    RECT 0 1124.375 0.070 1124.445 ;
    RECT 0 1124.515 0.070 1124.585 ;
    RECT 0 1124.655 0.070 1124.725 ;
    RECT 0 1124.795 0.070 1124.865 ;
    RECT 0 1124.935 0.070 1125.005 ;
    RECT 0 1125.075 0.070 1125.145 ;
    RECT 0 1125.215 0.070 1125.285 ;
    RECT 0 1125.355 0.070 1125.425 ;
    RECT 0 1125.495 0.070 1125.565 ;
    RECT 0 1125.635 0.070 1125.705 ;
    RECT 0 1125.775 0.070 1125.845 ;
    RECT 0 1125.915 0.070 1125.985 ;
    RECT 0 1126.055 0.070 1126.125 ;
    RECT 0 1126.195 0.070 1126.265 ;
    RECT 0 1126.335 0.070 1126.405 ;
    RECT 0 1126.475 0.070 1126.545 ;
    RECT 0 1126.615 0.070 1126.685 ;
    RECT 0 1126.755 0.070 1126.825 ;
    RECT 0 1126.895 0.070 1126.965 ;
    RECT 0 1127.035 0.070 1127.105 ;
    RECT 0 1127.175 0.070 1127.245 ;
    RECT 0 1127.315 0.070 1127.385 ;
    RECT 0 1127.455 0.070 1127.525 ;
    RECT 0 1127.595 0.070 1127.665 ;
    RECT 0 1127.735 0.070 1127.805 ;
    RECT 0 1127.875 0.070 1127.945 ;
    RECT 0 1128.015 0.070 1128.085 ;
    RECT 0 1128.155 0.070 1128.225 ;
    RECT 0 1128.295 0.070 1128.365 ;
    RECT 0 1128.435 0.070 1128.505 ;
    RECT 0 1128.575 0.070 1128.645 ;
    RECT 0 1128.715 0.070 1128.785 ;
    RECT 0 1128.855 0.070 1128.925 ;
    RECT 0 1128.995 0.070 1129.065 ;
    RECT 0 1129.135 0.070 1129.205 ;
    RECT 0 1129.275 0.070 1129.345 ;
    RECT 0 1129.415 0.070 1129.485 ;
    RECT 0 1129.555 0.070 1129.625 ;
    RECT 0 1129.695 0.070 1129.765 ;
    RECT 0 1129.835 0.070 1129.905 ;
    RECT 0 1129.975 0.070 1130.045 ;
    RECT 0 1130.115 0.070 1130.185 ;
    RECT 0 1130.255 0.070 1130.325 ;
    RECT 0 1130.395 0.070 1130.465 ;
    RECT 0 1130.535 0.070 1130.605 ;
    RECT 0 1130.675 0.070 1130.745 ;
    RECT 0 1130.815 0.070 1130.885 ;
    RECT 0 1130.955 0.070 1131.025 ;
    RECT 0 1131.095 0.070 1131.165 ;
    RECT 0 1131.235 0.070 1131.305 ;
    RECT 0 1131.375 0.070 1131.445 ;
    RECT 0 1131.515 0.070 1131.585 ;
    RECT 0 1131.655 0.070 1131.725 ;
    RECT 0 1131.795 0.070 1131.865 ;
    RECT 0 1131.935 0.070 1132.005 ;
    RECT 0 1132.075 0.070 1132.145 ;
    RECT 0 1132.215 0.070 1132.285 ;
    RECT 0 1132.355 0.070 1132.425 ;
    RECT 0 1132.495 0.070 1132.565 ;
    RECT 0 1132.635 0.070 1132.705 ;
    RECT 0 1132.775 0.070 1132.845 ;
    RECT 0 1132.915 0.070 1132.985 ;
    RECT 0 1133.055 0.070 1133.125 ;
    RECT 0 1133.195 0.070 1133.265 ;
    RECT 0 1133.335 0.070 1133.405 ;
    RECT 0 1133.475 0.070 1133.545 ;
    RECT 0 1133.615 0.070 1133.685 ;
    RECT 0 1133.755 0.070 1133.825 ;
    RECT 0 1133.895 0.070 1133.965 ;
    RECT 0 1134.035 0.070 1134.105 ;
    RECT 0 1134.175 0.070 1134.245 ;
    RECT 0 1134.315 0.070 1134.385 ;
    RECT 0 1134.455 0.070 1134.525 ;
    RECT 0 1134.595 0.070 1134.665 ;
    RECT 0 1134.735 0.070 1134.805 ;
    RECT 0 1134.875 0.070 1134.945 ;
    RECT 0 1135.015 0.070 1135.085 ;
    RECT 0 1135.155 0.070 1135.225 ;
    RECT 0 1135.295 0.070 1135.365 ;
    RECT 0 1135.435 0.070 1135.505 ;
    RECT 0 1135.575 0.070 1135.645 ;
    RECT 0 1135.715 0.070 1135.785 ;
    RECT 0 1135.855 0.070 1135.925 ;
    RECT 0 1135.995 0.070 1136.065 ;
    RECT 0 1136.135 0.070 1136.205 ;
    RECT 0 1136.275 0.070 1136.345 ;
    RECT 0 1136.415 0.070 1136.485 ;
    RECT 0 1136.555 0.070 1136.625 ;
    RECT 0 1136.695 0.070 1136.765 ;
    RECT 0 1136.835 0.070 1136.905 ;
    RECT 0 1136.975 0.070 1137.045 ;
    RECT 0 1137.115 0.070 1137.185 ;
    RECT 0 1137.255 0.070 1137.325 ;
    RECT 0 1137.395 0.070 1137.465 ;
    RECT 0 1137.535 0.070 1137.605 ;
    RECT 0 1137.675 0.070 1137.745 ;
    RECT 0 1137.815 0.070 1137.885 ;
    RECT 0 1137.955 0.070 1138.025 ;
    RECT 0 1138.095 0.070 1138.165 ;
    RECT 0 1138.235 0.070 1138.305 ;
    RECT 0 1138.375 0.070 1138.445 ;
    RECT 0 1138.515 0.070 1138.585 ;
    RECT 0 1138.655 0.070 1138.725 ;
    RECT 0 1138.795 0.070 1138.865 ;
    RECT 0 1138.935 0.070 1139.005 ;
    RECT 0 1139.075 0.070 1139.145 ;
    RECT 0 1139.215 0.070 1139.285 ;
    RECT 0 1139.355 0.070 1139.425 ;
    RECT 0 1139.495 0.070 1139.565 ;
    RECT 0 1139.635 0.070 1139.705 ;
    RECT 0 1139.775 0.070 1139.845 ;
    RECT 0 1139.915 0.070 1139.985 ;
    RECT 0 1140.055 0.070 1140.125 ;
    RECT 0 1140.195 0.070 1140.265 ;
    RECT 0 1140.335 0.070 1140.405 ;
    RECT 0 1140.475 0.070 1140.545 ;
    RECT 0 1140.615 0.070 1140.685 ;
    RECT 0 1140.755 0.070 1140.825 ;
    RECT 0 1140.895 0.070 1140.965 ;
    RECT 0 1141.035 0.070 1141.105 ;
    RECT 0 1141.175 0.070 1141.245 ;
    RECT 0 1141.315 0.070 1141.385 ;
    RECT 0 1141.455 0.070 1141.525 ;
    RECT 0 1141.595 0.070 1141.665 ;
    RECT 0 1141.735 0.070 1141.805 ;
    RECT 0 1141.875 0.070 1141.945 ;
    RECT 0 1142.015 0.070 1142.085 ;
    RECT 0 1142.155 0.070 1142.225 ;
    RECT 0 1142.295 0.070 1142.365 ;
    RECT 0 1142.435 0.070 1142.505 ;
    RECT 0 1142.575 0.070 1142.645 ;
    RECT 0 1142.715 0.070 1142.785 ;
    RECT 0 1142.855 0.070 1142.925 ;
    RECT 0 1142.995 0.070 1143.065 ;
    RECT 0 1143.135 0.070 1143.205 ;
    RECT 0 1143.275 0.070 1143.345 ;
    RECT 0 1143.415 0.070 1143.485 ;
    RECT 0 1143.555 0.070 1143.625 ;
    RECT 0 1143.695 0.070 1143.765 ;
    RECT 0 1143.835 0.070 1143.905 ;
    RECT 0 1143.975 0.070 1144.045 ;
    RECT 0 1144.115 0.070 1144.185 ;
    RECT 0 1144.255 0.070 1144.325 ;
    RECT 0 1144.395 0.070 1144.465 ;
    RECT 0 1144.535 0.070 1144.605 ;
    RECT 0 1144.675 0.070 1144.745 ;
    RECT 0 1144.815 0.070 1144.885 ;
    RECT 0 1144.955 0.070 1145.025 ;
    RECT 0 1145.095 0.070 1145.165 ;
    RECT 0 1145.235 0.070 1145.305 ;
    RECT 0 1145.375 0.070 1145.445 ;
    RECT 0 1145.515 0.070 1145.585 ;
    RECT 0 1145.655 0.070 1145.725 ;
    RECT 0 1145.795 0.070 1145.865 ;
    RECT 0 1145.935 0.070 1146.005 ;
    RECT 0 1146.075 0.070 1146.145 ;
    RECT 0 1146.215 0.070 1146.285 ;
    RECT 0 1146.355 0.070 1146.425 ;
    RECT 0 1146.495 0.070 1146.565 ;
    RECT 0 1146.635 0.070 1146.705 ;
    RECT 0 1146.775 0.070 1146.845 ;
    RECT 0 1146.915 0.070 1146.985 ;
    RECT 0 1147.055 0.070 1147.125 ;
    RECT 0 1147.195 0.070 1147.265 ;
    RECT 0 1147.335 0.070 1147.405 ;
    RECT 0 1147.475 0.070 1147.545 ;
    RECT 0 1147.615 0.070 1147.685 ;
    RECT 0 1147.755 0.070 1147.825 ;
    RECT 0 1147.895 0.070 1147.965 ;
    RECT 0 1148.035 0.070 1148.105 ;
    RECT 0 1148.175 0.070 1148.245 ;
    RECT 0 1148.315 0.070 1148.385 ;
    RECT 0 1148.455 0.070 1148.525 ;
    RECT 0 1148.595 0.070 1148.665 ;
    RECT 0 1148.735 0.070 1148.805 ;
    RECT 0 1148.875 0.070 1148.945 ;
    RECT 0 1149.015 0.070 1149.085 ;
    RECT 0 1149.155 0.070 1149.225 ;
    RECT 0 1149.295 0.070 1149.365 ;
    RECT 0 1149.435 0.070 1149.505 ;
    RECT 0 1149.575 0.070 1149.645 ;
    RECT 0 1149.715 0.070 1149.785 ;
    RECT 0 1149.855 0.070 1149.925 ;
    RECT 0 1149.995 0.070 1150.065 ;
    RECT 0 1150.135 0.070 1150.205 ;
    RECT 0 1150.275 0.070 1150.345 ;
    RECT 0 1150.415 0.070 1150.485 ;
    RECT 0 1150.555 0.070 1150.625 ;
    RECT 0 1150.695 0.070 1150.765 ;
    RECT 0 1150.835 0.070 1150.905 ;
    RECT 0 1150.975 0.070 1151.045 ;
    RECT 0 1151.115 0.070 1151.185 ;
    RECT 0 1151.255 0.070 1151.325 ;
    RECT 0 1151.395 0.070 1151.465 ;
    RECT 0 1151.535 0.070 1151.605 ;
    RECT 0 1151.675 0.070 1151.745 ;
    RECT 0 1151.815 0.070 1151.885 ;
    RECT 0 1151.955 0.070 1152.025 ;
    RECT 0 1152.095 0.070 1152.165 ;
    RECT 0 1152.235 0.070 1152.305 ;
    RECT 0 1152.375 0.070 1152.445 ;
    RECT 0 1152.515 0.070 1152.585 ;
    RECT 0 1152.655 0.070 1152.725 ;
    RECT 0 1152.795 0.070 1152.865 ;
    RECT 0 1152.935 0.070 1153.005 ;
    RECT 0 1153.075 0.070 1153.145 ;
    RECT 0 1153.215 0.070 1153.285 ;
    RECT 0 1153.355 0.070 1153.425 ;
    RECT 0 1153.495 0.070 1153.565 ;
    RECT 0 1153.635 0.070 1153.705 ;
    RECT 0 1153.775 0.070 1153.845 ;
    RECT 0 1153.915 0.070 1153.985 ;
    RECT 0 1154.055 0.070 1154.125 ;
    RECT 0 1154.195 0.070 1154.265 ;
    RECT 0 1154.335 0.070 1154.405 ;
    RECT 0 1154.475 0.070 1154.545 ;
    RECT 0 1154.615 0.070 1154.685 ;
    RECT 0 1154.755 0.070 1154.825 ;
    RECT 0 1154.895 0.070 1154.965 ;
    RECT 0 1155.035 0.070 1155.105 ;
    RECT 0 1155.175 0.070 1155.245 ;
    RECT 0 1155.315 0.070 1155.385 ;
    RECT 0 1155.455 0.070 1155.525 ;
    RECT 0 1155.595 0.070 1155.665 ;
    RECT 0 1155.735 0.070 1155.805 ;
    RECT 0 1155.875 0.070 1155.945 ;
    RECT 0 1156.015 0.070 1156.085 ;
    RECT 0 1156.155 0.070 1156.225 ;
    RECT 0 1156.295 0.070 1156.365 ;
    RECT 0 1156.435 0.070 1156.505 ;
    RECT 0 1156.575 0.070 1156.645 ;
    RECT 0 1156.715 0.070 1156.785 ;
    RECT 0 1156.855 0.070 1156.925 ;
    RECT 0 1156.995 0.070 1157.065 ;
    RECT 0 1157.135 0.070 1157.205 ;
    RECT 0 1157.275 0.070 1157.345 ;
    RECT 0 1157.415 0.070 1157.485 ;
    RECT 0 1157.555 0.070 1157.625 ;
    RECT 0 1157.695 0.070 1157.765 ;
    RECT 0 1157.835 0.070 1157.905 ;
    RECT 0 1157.975 0.070 1158.045 ;
    RECT 0 1158.115 0.070 1158.185 ;
    RECT 0 1158.255 0.070 1158.325 ;
    RECT 0 1158.395 0.070 1158.465 ;
    RECT 0 1158.535 0.070 1158.605 ;
    RECT 0 1158.675 0.070 1158.745 ;
    RECT 0 1158.815 0.070 1158.885 ;
    RECT 0 1158.955 0.070 1159.025 ;
    RECT 0 1159.095 0.070 1159.165 ;
    RECT 0 1159.235 0.070 1159.305 ;
    RECT 0 1159.375 0.070 1159.445 ;
    RECT 0 1159.515 0.070 1159.585 ;
    RECT 0 1159.655 0.070 1159.725 ;
    RECT 0 1159.795 0.070 1159.865 ;
    RECT 0 1159.935 0.070 1160.005 ;
    RECT 0 1160.075 0.070 1160.145 ;
    RECT 0 1160.215 0.070 1160.285 ;
    RECT 0 1160.355 0.070 1160.425 ;
    RECT 0 1160.495 0.070 1160.565 ;
    RECT 0 1160.635 0.070 1160.705 ;
    RECT 0 1160.775 0.070 1160.845 ;
    RECT 0 1160.915 0.070 1160.985 ;
    RECT 0 1161.055 0.070 1161.125 ;
    RECT 0 1161.195 0.070 1161.265 ;
    RECT 0 1161.335 0.070 1161.405 ;
    RECT 0 1161.475 0.070 1161.545 ;
    RECT 0 1161.615 0.070 1161.685 ;
    RECT 0 1161.755 0.070 1161.825 ;
    RECT 0 1161.895 0.070 1161.965 ;
    RECT 0 1162.035 0.070 1162.105 ;
    RECT 0 1162.175 0.070 1162.245 ;
    RECT 0 1162.315 0.070 1162.385 ;
    RECT 0 1162.455 0.070 1162.525 ;
    RECT 0 1162.595 0.070 1162.665 ;
    RECT 0 1162.735 0.070 1162.805 ;
    RECT 0 1162.875 0.070 1162.945 ;
    RECT 0 1163.015 0.070 1163.085 ;
    RECT 0 1163.155 0.070 1163.225 ;
    RECT 0 1163.295 0.070 1163.365 ;
    RECT 0 1163.435 0.070 1163.505 ;
    RECT 0 1163.575 0.070 1163.645 ;
    RECT 0 1163.715 0.070 1163.785 ;
    RECT 0 1163.855 0.070 1163.925 ;
    RECT 0 1163.995 0.070 1164.065 ;
    RECT 0 1164.135 0.070 1164.205 ;
    RECT 0 1164.275 0.070 1164.345 ;
    RECT 0 1164.415 0.070 1164.485 ;
    RECT 0 1164.555 0.070 1164.625 ;
    RECT 0 1164.695 0.070 1164.765 ;
    RECT 0 1164.835 0.070 1164.905 ;
    RECT 0 1164.975 0.070 1165.045 ;
    RECT 0 1165.115 0.070 1165.185 ;
    RECT 0 1165.255 0.070 1165.325 ;
    RECT 0 1165.395 0.070 1165.465 ;
    RECT 0 1165.535 0.070 1165.605 ;
    RECT 0 1165.675 0.070 1165.745 ;
    RECT 0 1165.815 0.070 1165.885 ;
    RECT 0 1165.955 0.070 1166.025 ;
    RECT 0 1166.095 0.070 1166.165 ;
    RECT 0 1166.235 0.070 1166.305 ;
    RECT 0 1166.375 0.070 1166.445 ;
    RECT 0 1166.515 0.070 1166.585 ;
    RECT 0 1166.655 0.070 1166.725 ;
    RECT 0 1166.795 0.070 1166.865 ;
    RECT 0 1166.935 0.070 1167.005 ;
    RECT 0 1167.075 0.070 1167.145 ;
    RECT 0 1167.215 0.070 1167.285 ;
    RECT 0 1167.355 0.070 1167.425 ;
    RECT 0 1167.495 0.070 1167.565 ;
    RECT 0 1167.635 0.070 1167.705 ;
    RECT 0 1167.775 0.070 1167.845 ;
    RECT 0 1167.915 0.070 1167.985 ;
    RECT 0 1168.055 0.070 1168.125 ;
    RECT 0 1168.195 0.070 1168.265 ;
    RECT 0 1168.335 0.070 1168.405 ;
    RECT 0 1168.475 0.070 1168.545 ;
    RECT 0 1168.615 0.070 1168.685 ;
    RECT 0 1168.755 0.070 1168.825 ;
    RECT 0 1168.895 0.070 1168.965 ;
    RECT 0 1169.035 0.070 1169.105 ;
    RECT 0 1169.175 0.070 1169.245 ;
    RECT 0 1169.315 0.070 1169.385 ;
    RECT 0 1169.455 0.070 1169.525 ;
    RECT 0 1169.595 0.070 1169.665 ;
    RECT 0 1169.735 0.070 1169.805 ;
    RECT 0 1169.875 0.070 1169.945 ;
    RECT 0 1170.015 0.070 1170.085 ;
    RECT 0 1170.155 0.070 1170.225 ;
    RECT 0 1170.295 0.070 1170.365 ;
    RECT 0 1170.435 0.070 1170.505 ;
    RECT 0 1170.575 0.070 1170.645 ;
    RECT 0 1170.715 0.070 1170.785 ;
    RECT 0 1170.855 0.070 1170.925 ;
    RECT 0 1170.995 0.070 1171.065 ;
    RECT 0 1171.135 0.070 1171.205 ;
    RECT 0 1171.275 0.070 1171.345 ;
    RECT 0 1171.415 0.070 1171.485 ;
    RECT 0 1171.555 0.070 1171.625 ;
    RECT 0 1171.695 0.070 1171.765 ;
    RECT 0 1171.835 0.070 1171.905 ;
    RECT 0 1171.975 0.070 1172.045 ;
    RECT 0 1172.115 0.070 1172.185 ;
    RECT 0 1172.255 0.070 1172.325 ;
    RECT 0 1172.395 0.070 1172.465 ;
    RECT 0 1172.535 0.070 1172.605 ;
    RECT 0 1172.675 0.070 1172.745 ;
    RECT 0 1172.815 0.070 1172.885 ;
    RECT 0 1172.955 0.070 1173.025 ;
    RECT 0 1173.095 0.070 1173.165 ;
    RECT 0 1173.235 0.070 1173.305 ;
    RECT 0 1173.375 0.070 1173.445 ;
    RECT 0 1173.515 0.070 1173.585 ;
    RECT 0 1173.655 0.070 1173.725 ;
    RECT 0 1173.795 0.070 1173.865 ;
    RECT 0 1173.935 0.070 1174.005 ;
    RECT 0 1174.075 0.070 1174.145 ;
    RECT 0 1174.215 0.070 1174.285 ;
    RECT 0 1174.355 0.070 1174.425 ;
    RECT 0 1174.495 0.070 1174.565 ;
    RECT 0 1174.635 0.070 1174.705 ;
    RECT 0 1174.775 0.070 1174.845 ;
    RECT 0 1174.915 0.070 1174.985 ;
    RECT 0 1175.055 0.070 1175.125 ;
    RECT 0 1175.195 0.070 1175.265 ;
    RECT 0 1175.335 0.070 1175.405 ;
    RECT 0 1175.475 0.070 1175.545 ;
    RECT 0 1175.615 0.070 1175.685 ;
    RECT 0 1175.755 0.070 1175.825 ;
    RECT 0 1175.895 0.070 1175.965 ;
    RECT 0 1176.035 0.070 1176.105 ;
    RECT 0 1176.175 0.070 1176.245 ;
    RECT 0 1176.315 0.070 1176.385 ;
    RECT 0 1176.455 0.070 1176.525 ;
    RECT 0 1176.595 0.070 1176.665 ;
    RECT 0 1176.735 0.070 1176.805 ;
    RECT 0 1176.875 0.070 1176.945 ;
    RECT 0 1177.015 0.070 1177.085 ;
    RECT 0 1177.155 0.070 1177.225 ;
    RECT 0 1177.295 0.070 1177.365 ;
    RECT 0 1177.435 0.070 1177.505 ;
    RECT 0 1177.575 0.070 1177.645 ;
    RECT 0 1177.715 0.070 1177.785 ;
    RECT 0 1177.855 0.070 1177.925 ;
    RECT 0 1177.995 0.070 1178.065 ;
    RECT 0 1178.135 0.070 1178.205 ;
    RECT 0 1178.275 0.070 1178.345 ;
    RECT 0 1178.415 0.070 1178.485 ;
    RECT 0 1178.555 0.070 1178.625 ;
    RECT 0 1178.695 0.070 1178.765 ;
    RECT 0 1178.835 0.070 1178.905 ;
    RECT 0 1178.975 0.070 1179.045 ;
    RECT 0 1179.115 0.070 1179.185 ;
    RECT 0 1179.255 0.070 1179.325 ;
    RECT 0 1179.395 0.070 1179.465 ;
    RECT 0 1179.535 0.070 1179.605 ;
    RECT 0 1179.675 0.070 1179.745 ;
    RECT 0 1179.815 0.070 1179.885 ;
    RECT 0 1179.955 0.070 1180.025 ;
    RECT 0 1180.095 0.070 1180.165 ;
    RECT 0 1180.235 0.070 1180.305 ;
    RECT 0 1180.375 0.070 1180.445 ;
    RECT 0 1180.515 0.070 1180.585 ;
    RECT 0 1180.655 0.070 1180.725 ;
    RECT 0 1180.795 0.070 1180.865 ;
    RECT 0 1180.935 0.070 1181.005 ;
    RECT 0 1181.075 0.070 1181.145 ;
    RECT 0 1181.215 0.070 1181.285 ;
    RECT 0 1181.355 0.070 1181.425 ;
    RECT 0 1181.495 0.070 1181.565 ;
    RECT 0 1181.635 0.070 1181.705 ;
    RECT 0 1181.775 0.070 1181.845 ;
    RECT 0 1181.915 0.070 1181.985 ;
    RECT 0 1182.055 0.070 1182.125 ;
    RECT 0 1182.195 0.070 1182.265 ;
    RECT 0 1182.335 0.070 1182.405 ;
    RECT 0 1182.475 0.070 1182.545 ;
    RECT 0 1182.615 0.070 1182.685 ;
    RECT 0 1182.755 0.070 1182.825 ;
    RECT 0 1182.895 0.070 1182.965 ;
    RECT 0 1183.035 0.070 1183.105 ;
    RECT 0 1183.175 0.070 1183.245 ;
    RECT 0 1183.315 0.070 1183.385 ;
    RECT 0 1183.455 0.070 1183.525 ;
    RECT 0 1183.595 0.070 1183.665 ;
    RECT 0 1183.735 0.070 1183.805 ;
    RECT 0 1183.875 0.070 1183.945 ;
    RECT 0 1184.015 0.070 1184.085 ;
    RECT 0 1184.155 0.070 1184.225 ;
    RECT 0 1184.295 0.070 1184.365 ;
    RECT 0 1184.435 0.070 1184.505 ;
    RECT 0 1184.575 0.070 1184.645 ;
    RECT 0 1184.715 0.070 1184.785 ;
    RECT 0 1184.855 0.070 1184.925 ;
    RECT 0 1184.995 0.070 1185.065 ;
    RECT 0 1185.135 0.070 1185.205 ;
    RECT 0 1185.275 0.070 1185.345 ;
    RECT 0 1185.415 0.070 1185.485 ;
    RECT 0 1185.555 0.070 1185.625 ;
    RECT 0 1185.695 0.070 1185.765 ;
    RECT 0 1185.835 0.070 1185.905 ;
    RECT 0 1185.975 0.070 1186.045 ;
    RECT 0 1186.115 0.070 1186.185 ;
    RECT 0 1186.255 0.070 1186.325 ;
    RECT 0 1186.395 0.070 1186.465 ;
    RECT 0 1186.535 0.070 1186.605 ;
    RECT 0 1186.675 0.070 1186.745 ;
    RECT 0 1186.815 0.070 1186.885 ;
    RECT 0 1186.955 0.070 1187.025 ;
    RECT 0 1187.095 0.070 1187.165 ;
    RECT 0 1187.235 0.070 1187.305 ;
    RECT 0 1187.375 0.070 1187.445 ;
    RECT 0 1187.515 0.070 1187.585 ;
    RECT 0 1187.655 0.070 1187.725 ;
    RECT 0 1187.795 0.070 1187.865 ;
    RECT 0 1187.935 0.070 1188.005 ;
    RECT 0 1188.075 0.070 1188.145 ;
    RECT 0 1188.215 0.070 1188.285 ;
    RECT 0 1188.355 0.070 1188.425 ;
    RECT 0 1188.495 0.070 1188.565 ;
    RECT 0 1188.635 0.070 1188.705 ;
    RECT 0 1188.775 0.070 1188.845 ;
    RECT 0 1188.915 0.070 1188.985 ;
    RECT 0 1189.055 0.070 1189.125 ;
    RECT 0 1189.195 0.070 1189.265 ;
    RECT 0 1189.335 0.070 1189.405 ;
    RECT 0 1189.475 0.070 1189.545 ;
    RECT 0 1189.615 0.070 1189.685 ;
    RECT 0 1189.755 0.070 1189.825 ;
    RECT 0 1189.895 0.070 1189.965 ;
    RECT 0 1190.035 0.070 1190.105 ;
    RECT 0 1190.175 0.070 1190.245 ;
    RECT 0 1190.315 0.070 1190.385 ;
    RECT 0 1190.455 0.070 1190.525 ;
    RECT 0 1190.595 0.070 1190.665 ;
    RECT 0 1190.735 0.070 1190.805 ;
    RECT 0 1190.875 0.070 1190.945 ;
    RECT 0 1191.015 0.070 1191.085 ;
    RECT 0 1191.155 0.070 1191.225 ;
    RECT 0 1191.295 0.070 1191.365 ;
    RECT 0 1191.435 0.070 1191.505 ;
    RECT 0 1191.575 0.070 1191.645 ;
    RECT 0 1191.715 0.070 1191.785 ;
    RECT 0 1191.855 0.070 1191.925 ;
    RECT 0 1191.995 0.070 1192.065 ;
    RECT 0 1192.135 0.070 1192.205 ;
    RECT 0 1192.275 0.070 1192.345 ;
    RECT 0 1192.415 0.070 1192.485 ;
    RECT 0 1192.555 0.070 1192.625 ;
    RECT 0 1192.695 0.070 1192.765 ;
    RECT 0 1192.835 0.070 1192.905 ;
    RECT 0 1192.975 0.070 1193.045 ;
    RECT 0 1193.115 0.070 1193.185 ;
    RECT 0 1193.255 0.070 1193.325 ;
    RECT 0 1193.395 0.070 1193.465 ;
    RECT 0 1193.535 0.070 1193.605 ;
    RECT 0 1193.675 0.070 1193.745 ;
    RECT 0 1193.815 0.070 1193.885 ;
    RECT 0 1193.955 0.070 1194.025 ;
    RECT 0 1194.095 0.070 1194.165 ;
    RECT 0 1194.235 0.070 1194.305 ;
    RECT 0 1194.375 0.070 1194.445 ;
    RECT 0 1194.515 0.070 1194.585 ;
    RECT 0 1194.655 0.070 1194.725 ;
    RECT 0 1194.795 0.070 1194.865 ;
    RECT 0 1194.935 0.070 1195.005 ;
    RECT 0 1195.075 0.070 1195.145 ;
    RECT 0 1195.215 0.070 1195.285 ;
    RECT 0 1195.355 0.070 1195.425 ;
    RECT 0 1195.495 0.070 1195.565 ;
    RECT 0 1195.635 0.070 1195.705 ;
    RECT 0 1195.775 0.070 1195.845 ;
    RECT 0 1195.915 0.070 1195.985 ;
    RECT 0 1196.055 0.070 1196.125 ;
    RECT 0 1196.195 0.070 1196.265 ;
    RECT 0 1196.335 0.070 1196.405 ;
    RECT 0 1196.475 0.070 1196.545 ;
    RECT 0 1196.615 0.070 1196.685 ;
    RECT 0 1196.755 0.070 1196.825 ;
    RECT 0 1196.895 0.070 1196.965 ;
    RECT 0 1197.035 0.070 1197.105 ;
    RECT 0 1197.175 0.070 1197.245 ;
    RECT 0 1197.315 0.070 1197.385 ;
    RECT 0 1197.455 0.070 1197.525 ;
    RECT 0 1197.595 0.070 1197.665 ;
    RECT 0 1197.735 0.070 1197.805 ;
    RECT 0 1197.875 0.070 1197.945 ;
    RECT 0 1198.015 0.070 1198.085 ;
    RECT 0 1198.155 0.070 1198.225 ;
    RECT 0 1198.295 0.070 1198.365 ;
    RECT 0 1198.435 0.070 1198.505 ;
    RECT 0 1198.575 0.070 1198.645 ;
    RECT 0 1198.715 0.070 1198.785 ;
    RECT 0 1198.855 0.070 1198.925 ;
    RECT 0 1198.995 0.070 1199.065 ;
    RECT 0 1199.135 0.070 1199.205 ;
    RECT 0 1199.275 0.070 1199.345 ;
    RECT 0 1199.415 0.070 1199.485 ;
    RECT 0 1199.555 0.070 1199.625 ;
    RECT 0 1199.695 0.070 1199.765 ;
    RECT 0 1199.835 0.070 1199.905 ;
    RECT 0 1199.975 0.070 1200.045 ;
    RECT 0 1200.115 0.070 1200.185 ;
    RECT 0 1200.255 0.070 1200.325 ;
    RECT 0 1200.395 0.070 1200.465 ;
    RECT 0 1200.535 0.070 1200.605 ;
    RECT 0 1200.675 0.070 1200.745 ;
    RECT 0 1200.815 0.070 1200.885 ;
    RECT 0 1200.955 0.070 1201.025 ;
    RECT 0 1201.095 0.070 1201.165 ;
    RECT 0 1201.235 0.070 1201.305 ;
    RECT 0 1201.375 0.070 1201.445 ;
    RECT 0 1201.515 0.070 1201.585 ;
    RECT 0 1201.655 0.070 1201.725 ;
    RECT 0 1201.795 0.070 1201.865 ;
    RECT 0 1201.935 0.070 1202.005 ;
    RECT 0 1202.075 0.070 1202.145 ;
    RECT 0 1202.215 0.070 1202.285 ;
    RECT 0 1202.355 0.070 1202.425 ;
    RECT 0 1202.495 0.070 1202.565 ;
    RECT 0 1202.635 0.070 1202.705 ;
    RECT 0 1202.775 0.070 1202.845 ;
    RECT 0 1202.915 0.070 1202.985 ;
    RECT 0 1203.055 0.070 1203.125 ;
    RECT 0 1203.195 0.070 1203.265 ;
    RECT 0 1203.335 0.070 1203.405 ;
    RECT 0 1203.475 0.070 1203.545 ;
    RECT 0 1203.615 0.070 1203.685 ;
    RECT 0 1203.755 0.070 1203.825 ;
    RECT 0 1203.895 0.070 1203.965 ;
    RECT 0 1204.035 0.070 1204.105 ;
    RECT 0 1204.175 0.070 1204.245 ;
    RECT 0 1204.315 0.070 1204.385 ;
    RECT 0 1204.455 0.070 1204.525 ;
    RECT 0 1204.595 0.070 1204.665 ;
    RECT 0 1204.735 0.070 1204.805 ;
    RECT 0 1204.875 0.070 1204.945 ;
    RECT 0 1205.015 0.070 1205.085 ;
    RECT 0 1205.155 0.070 1205.225 ;
    RECT 0 1205.295 0.070 1205.365 ;
    RECT 0 1205.435 0.070 1205.505 ;
    RECT 0 1205.575 0.070 1205.645 ;
    RECT 0 1205.715 0.070 1205.785 ;
    RECT 0 1205.855 0.070 1205.925 ;
    RECT 0 1205.995 0.070 1206.065 ;
    RECT 0 1206.135 0.070 1206.205 ;
    RECT 0 1206.275 0.070 1206.345 ;
    RECT 0 1206.415 0.070 1206.485 ;
    RECT 0 1206.555 0.070 1206.625 ;
    RECT 0 1206.695 0.070 1206.765 ;
    RECT 0 1206.835 0.070 1206.905 ;
    RECT 0 1206.975 0.070 1207.045 ;
    RECT 0 1207.115 0.070 1207.185 ;
    RECT 0 1207.255 0.070 1207.325 ;
    RECT 0 1207.395 0.070 1207.465 ;
    RECT 0 1207.535 0.070 1207.605 ;
    RECT 0 1207.675 0.070 1207.745 ;
    RECT 0 1207.815 0.070 1207.885 ;
    RECT 0 1207.955 0.070 1208.025 ;
    RECT 0 1208.095 0.070 1208.165 ;
    RECT 0 1208.235 0.070 1208.305 ;
    RECT 0 1208.375 0.070 1208.445 ;
    RECT 0 1208.515 0.070 1208.585 ;
    RECT 0 1208.655 0.070 1208.725 ;
    RECT 0 1208.795 0.070 1208.865 ;
    RECT 0 1208.935 0.070 1209.005 ;
    RECT 0 1209.075 0.070 1209.145 ;
    RECT 0 1209.215 0.070 1209.285 ;
    RECT 0 1209.355 0.070 1209.425 ;
    RECT 0 1209.495 0.070 1209.565 ;
    RECT 0 1209.635 0.070 1209.705 ;
    RECT 0 1209.775 0.070 1209.845 ;
    RECT 0 1209.915 0.070 1209.985 ;
    RECT 0 1210.055 0.070 1210.125 ;
    RECT 0 1210.195 0.070 1210.265 ;
    RECT 0 1210.335 0.070 1210.405 ;
    RECT 0 1210.475 0.070 1210.545 ;
    RECT 0 1210.615 0.070 1210.685 ;
    RECT 0 1210.755 0.070 1210.825 ;
    RECT 0 1210.895 0.070 1210.965 ;
    RECT 0 1211.035 0.070 1211.105 ;
    RECT 0 1211.175 0.070 1211.245 ;
    RECT 0 1211.315 0.070 1211.385 ;
    RECT 0 1211.455 0.070 1211.525 ;
    RECT 0 1211.595 0.070 1211.665 ;
    RECT 0 1211.735 0.070 1211.805 ;
    RECT 0 1211.875 0.070 1211.945 ;
    RECT 0 1212.015 0.070 1212.085 ;
    RECT 0 1212.155 0.070 1212.225 ;
    RECT 0 1212.295 0.070 1212.365 ;
    RECT 0 1212.435 0.070 1212.505 ;
    RECT 0 1212.575 0.070 1212.645 ;
    RECT 0 1212.715 0.070 1212.785 ;
    RECT 0 1212.855 0.070 1212.925 ;
    RECT 0 1212.995 0.070 1213.065 ;
    RECT 0 1213.135 0.070 1213.205 ;
    RECT 0 1213.275 0.070 1213.345 ;
    RECT 0 1213.415 0.070 1213.485 ;
    RECT 0 1213.555 0.070 1213.625 ;
    RECT 0 1213.695 0.070 1213.765 ;
    RECT 0 1213.835 0.070 1213.905 ;
    RECT 0 1213.975 0.070 1214.045 ;
    RECT 0 1214.115 0.070 1214.185 ;
    RECT 0 1214.255 0.070 1214.325 ;
    RECT 0 1214.395 0.070 1214.465 ;
    RECT 0 1214.535 0.070 1214.605 ;
    RECT 0 1214.675 0.070 1214.745 ;
    RECT 0 1214.815 0.070 1214.885 ;
    RECT 0 1214.955 0.070 1215.025 ;
    RECT 0 1215.095 0.070 1215.165 ;
    RECT 0 1215.235 0.070 1215.305 ;
    RECT 0 1215.375 0.070 1215.445 ;
    RECT 0 1215.515 0.070 1215.585 ;
    RECT 0 1215.655 0.070 1215.725 ;
    RECT 0 1215.795 0.070 1215.865 ;
    RECT 0 1215.935 0.070 1216.005 ;
    RECT 0 1216.075 0.070 1216.145 ;
    RECT 0 1216.215 0.070 1216.285 ;
    RECT 0 1216.355 0.070 1216.425 ;
    RECT 0 1216.495 0.070 1216.565 ;
    RECT 0 1216.635 0.070 1216.705 ;
    RECT 0 1216.775 0.070 1216.845 ;
    RECT 0 1216.915 0.070 1216.985 ;
    RECT 0 1217.055 0.070 1217.125 ;
    RECT 0 1217.195 0.070 1217.265 ;
    RECT 0 1217.335 0.070 1217.405 ;
    RECT 0 1217.475 0.070 1217.545 ;
    RECT 0 1217.615 0.070 1217.685 ;
    RECT 0 1217.755 0.070 1217.825 ;
    RECT 0 1217.895 0.070 1217.965 ;
    RECT 0 1218.035 0.070 1218.105 ;
    RECT 0 1218.175 0.070 1218.245 ;
    RECT 0 1218.315 0.070 1218.385 ;
    RECT 0 1218.455 0.070 1218.525 ;
    RECT 0 1218.595 0.070 1218.665 ;
    RECT 0 1218.735 0.070 1218.805 ;
    RECT 0 1218.875 0.070 1218.945 ;
    RECT 0 1219.015 0.070 1219.085 ;
    RECT 0 1219.155 0.070 1219.225 ;
    RECT 0 1219.295 0.070 1219.365 ;
    RECT 0 1219.435 0.070 1219.505 ;
    RECT 0 1219.575 0.070 1219.645 ;
    RECT 0 1219.715 0.070 1219.785 ;
    RECT 0 1219.855 0.070 1219.925 ;
    RECT 0 1219.995 0.070 1220.065 ;
    RECT 0 1220.135 0.070 1220.205 ;
    RECT 0 1220.275 0.070 1220.345 ;
    RECT 0 1220.415 0.070 1220.485 ;
    RECT 0 1220.555 0.070 1220.625 ;
    RECT 0 1220.695 0.070 1220.765 ;
    RECT 0 1220.835 0.070 1220.905 ;
    RECT 0 1220.975 0.070 1221.045 ;
    RECT 0 1221.115 0.070 1221.185 ;
    RECT 0 1221.255 0.070 1221.325 ;
    RECT 0 1221.395 0.070 1221.465 ;
    RECT 0 1221.535 0.070 1221.605 ;
    RECT 0 1221.675 0.070 1221.745 ;
    RECT 0 1221.815 0.070 1221.885 ;
    RECT 0 1221.955 0.070 1222.025 ;
    RECT 0 1222.095 0.070 1222.165 ;
    RECT 0 1222.235 0.070 1222.305 ;
    RECT 0 1222.375 0.070 1222.445 ;
    RECT 0 1222.515 0.070 1222.585 ;
    RECT 0 1222.655 0.070 1222.725 ;
    RECT 0 1222.795 0.070 1222.865 ;
    RECT 0 1222.935 0.070 1223.005 ;
    RECT 0 1223.075 0.070 1223.145 ;
    RECT 0 1223.215 0.070 1223.285 ;
    RECT 0 1223.355 0.070 1223.425 ;
    RECT 0 1223.495 0.070 1223.565 ;
    RECT 0 1223.635 0.070 1223.705 ;
    RECT 0 1223.775 0.070 1223.845 ;
    RECT 0 1223.915 0.070 1223.985 ;
    RECT 0 1224.055 0.070 1224.125 ;
    RECT 0 1224.195 0.070 1224.265 ;
    RECT 0 1224.335 0.070 1224.405 ;
    RECT 0 1224.475 0.070 1224.545 ;
    RECT 0 1224.615 0.070 1224.685 ;
    RECT 0 1224.755 0.070 1224.825 ;
    RECT 0 1224.895 0.070 1224.965 ;
    RECT 0 1225.035 0.070 1225.105 ;
    RECT 0 1225.175 0.070 1225.245 ;
    RECT 0 1225.315 0.070 1225.385 ;
    RECT 0 1225.455 0.070 1225.525 ;
    RECT 0 1225.595 0.070 1225.665 ;
    RECT 0 1225.735 0.070 1225.805 ;
    RECT 0 1225.875 0.070 1225.945 ;
    RECT 0 1226.015 0.070 1226.085 ;
    RECT 0 1226.155 0.070 1226.225 ;
    RECT 0 1226.295 0.070 1226.365 ;
    RECT 0 1226.435 0.070 1226.505 ;
    RECT 0 1226.575 0.070 1226.645 ;
    RECT 0 1226.715 0.070 1226.785 ;
    RECT 0 1226.855 0.070 1226.925 ;
    RECT 0 1226.995 0.070 1227.065 ;
    RECT 0 1227.135 0.070 1227.205 ;
    RECT 0 1227.275 0.070 1227.345 ;
    RECT 0 1227.415 0.070 1227.485 ;
    RECT 0 1227.555 0.070 1227.625 ;
    RECT 0 1227.695 0.070 1227.765 ;
    RECT 0 1227.835 0.070 1227.905 ;
    RECT 0 1227.975 0.070 1228.045 ;
    RECT 0 1228.115 0.070 1228.185 ;
    RECT 0 1228.255 0.070 1228.325 ;
    RECT 0 1228.395 0.070 1228.465 ;
    RECT 0 1228.535 0.070 1228.605 ;
    RECT 0 1228.675 0.070 1228.745 ;
    RECT 0 1228.815 0.070 1228.885 ;
    RECT 0 1228.955 0.070 1229.025 ;
    RECT 0 1229.095 0.070 1229.165 ;
    RECT 0 1229.235 0.070 1229.305 ;
    RECT 0 1229.375 0.070 1229.445 ;
    RECT 0 1229.515 0.070 1229.585 ;
    RECT 0 1229.655 0.070 1229.725 ;
    RECT 0 1229.795 0.070 1229.865 ;
    RECT 0 1229.935 0.070 1230.005 ;
    RECT 0 1230.075 0.070 1230.145 ;
    RECT 0 1230.215 0.070 1230.285 ;
    RECT 0 1230.355 0.070 1230.425 ;
    RECT 0 1230.495 0.070 1230.565 ;
    RECT 0 1230.635 0.070 1230.705 ;
    RECT 0 1230.775 0.070 1230.845 ;
    RECT 0 1230.915 0.070 1230.985 ;
    RECT 0 1231.055 0.070 1231.125 ;
    RECT 0 1231.195 0.070 1231.265 ;
    RECT 0 1231.335 0.070 1231.405 ;
    RECT 0 1231.475 0.070 1231.545 ;
    RECT 0 1231.615 0.070 1231.685 ;
    RECT 0 1231.755 0.070 1231.825 ;
    RECT 0 1231.895 0.070 1231.965 ;
    RECT 0 1232.035 0.070 1232.105 ;
    RECT 0 1232.175 0.070 1232.245 ;
    RECT 0 1232.315 0.070 1232.385 ;
    RECT 0 1232.455 0.070 1232.525 ;
    RECT 0 1232.595 0.070 1232.665 ;
    RECT 0 1232.735 0.070 1232.805 ;
    RECT 0 1232.875 0.070 1232.945 ;
    RECT 0 1233.015 0.070 1233.085 ;
    RECT 0 1233.155 0.070 1233.225 ;
    RECT 0 1233.295 0.070 1233.365 ;
    RECT 0 1233.435 0.070 1233.505 ;
    RECT 0 1233.575 0.070 1233.645 ;
    RECT 0 1233.715 0.070 1233.785 ;
    RECT 0 1233.855 0.070 1233.925 ;
    RECT 0 1233.995 0.070 1234.065 ;
    RECT 0 1234.135 0.070 1234.205 ;
    RECT 0 1234.275 0.070 1234.345 ;
    RECT 0 1234.415 0.070 1234.485 ;
    RECT 0 1234.555 0.070 1234.625 ;
    RECT 0 1234.695 0.070 1234.765 ;
    RECT 0 1234.835 0.070 1234.905 ;
    RECT 0 1234.975 0.070 1235.045 ;
    RECT 0 1235.115 0.070 1235.185 ;
    RECT 0 1235.255 0.070 1235.325 ;
    RECT 0 1235.395 0.070 1235.465 ;
    RECT 0 1235.535 0.070 1235.605 ;
    RECT 0 1235.675 0.070 1235.745 ;
    RECT 0 1235.815 0.070 1235.885 ;
    RECT 0 1235.955 0.070 1236.025 ;
    RECT 0 1236.095 0.070 1236.165 ;
    RECT 0 1236.235 0.070 1236.305 ;
    RECT 0 1236.375 0.070 1236.445 ;
    RECT 0 1236.515 0.070 1236.585 ;
    RECT 0 1236.655 0.070 1236.725 ;
    RECT 0 1236.795 0.070 1236.865 ;
    RECT 0 1236.935 0.070 1237.005 ;
    RECT 0 1237.075 0.070 1237.145 ;
    RECT 0 1237.215 0.070 1237.285 ;
    RECT 0 1237.355 0.070 1237.425 ;
    RECT 0 1237.495 0.070 1237.565 ;
    RECT 0 1237.635 0.070 1237.705 ;
    RECT 0 1237.775 0.070 1237.845 ;
    RECT 0 1237.915 0.070 1237.985 ;
    RECT 0 1238.055 0.070 1238.125 ;
    RECT 0 1238.195 0.070 1238.265 ;
    RECT 0 1238.335 0.070 1238.405 ;
    RECT 0 1238.475 0.070 1238.545 ;
    RECT 0 1238.615 0.070 1238.685 ;
    RECT 0 1238.755 0.070 1238.825 ;
    RECT 0 1238.895 0.070 1238.965 ;
    RECT 0 1239.035 0.070 1239.105 ;
    RECT 0 1239.175 0.070 1239.245 ;
    RECT 0 1239.315 0.070 1239.385 ;
    RECT 0 1239.455 0.070 1239.525 ;
    RECT 0 1239.595 0.070 1239.665 ;
    RECT 0 1239.735 0.070 1239.805 ;
    RECT 0 1239.875 0.070 1239.945 ;
    RECT 0 1240.015 0.070 1240.085 ;
    RECT 0 1240.155 0.070 1240.225 ;
    RECT 0 1240.295 0.070 1240.365 ;
    RECT 0 1240.435 0.070 1240.505 ;
    RECT 0 1240.575 0.070 1240.645 ;
    RECT 0 1240.715 0.070 1240.785 ;
    RECT 0 1240.855 0.070 1240.925 ;
    RECT 0 1240.995 0.070 1241.065 ;
    RECT 0 1241.135 0.070 1241.205 ;
    RECT 0 1241.275 0.070 1241.345 ;
    RECT 0 1241.415 0.070 1241.485 ;
    RECT 0 1241.555 0.070 1241.625 ;
    RECT 0 1241.695 0.070 1241.765 ;
    RECT 0 1241.835 0.070 1241.905 ;
    RECT 0 1241.975 0.070 1242.045 ;
    RECT 0 1242.115 0.070 1242.185 ;
    RECT 0 1242.255 0.070 1242.325 ;
    RECT 0 1242.395 0.070 1242.465 ;
    RECT 0 1242.535 0.070 1242.605 ;
    RECT 0 1242.675 0.070 1242.745 ;
    RECT 0 1242.815 0.070 1242.885 ;
    RECT 0 1242.955 0.070 1243.025 ;
    RECT 0 1243.095 0.070 1243.165 ;
    RECT 0 1243.235 0.070 1243.305 ;
    RECT 0 1243.375 0.070 1243.445 ;
    RECT 0 1243.515 0.070 1243.585 ;
    RECT 0 1243.655 0.070 1243.725 ;
    RECT 0 1243.795 0.070 1243.865 ;
    RECT 0 1243.935 0.070 1244.005 ;
    RECT 0 1244.075 0.070 1244.145 ;
    RECT 0 1244.215 0.070 1244.285 ;
    RECT 0 1244.355 0.070 1244.425 ;
    RECT 0 1244.495 0.070 1244.565 ;
    RECT 0 1244.635 0.070 1244.705 ;
    RECT 0 1244.775 0.070 1244.845 ;
    RECT 0 1244.915 0.070 1244.985 ;
    RECT 0 1245.055 0.070 1245.125 ;
    RECT 0 1245.195 0.070 1245.265 ;
    RECT 0 1245.335 0.070 1245.405 ;
    RECT 0 1245.475 0.070 1245.545 ;
    RECT 0 1245.615 0.070 1245.685 ;
    RECT 0 1245.755 0.070 1245.825 ;
    RECT 0 1245.895 0.070 1245.965 ;
    RECT 0 1246.035 0.070 1246.105 ;
    RECT 0 1246.175 0.070 1246.245 ;
    RECT 0 1246.315 0.070 1246.385 ;
    RECT 0 1246.455 0.070 1246.525 ;
    RECT 0 1246.595 0.070 1246.665 ;
    RECT 0 1246.735 0.070 1246.805 ;
    RECT 0 1246.875 0.070 1246.945 ;
    RECT 0 1247.015 0.070 1247.085 ;
    RECT 0 1247.155 0.070 1247.225 ;
    RECT 0 1247.295 0.070 1247.365 ;
    RECT 0 1247.435 0.070 1247.505 ;
    RECT 0 1247.575 0.070 1247.645 ;
    RECT 0 1247.715 0.070 1247.785 ;
    RECT 0 1247.855 0.070 1247.925 ;
    RECT 0 1247.995 0.070 1248.065 ;
    RECT 0 1248.135 0.070 1248.205 ;
    RECT 0 1248.275 0.070 1248.345 ;
    RECT 0 1248.415 0.070 1248.485 ;
    RECT 0 1248.555 0.070 1248.625 ;
    RECT 0 1248.695 0.070 1248.765 ;
    RECT 0 1248.835 0.070 1248.905 ;
    RECT 0 1248.975 0.070 1249.045 ;
    RECT 0 1249.115 0.070 1249.185 ;
    RECT 0 1249.255 0.070 1249.325 ;
    RECT 0 1249.395 0.070 1249.465 ;
    RECT 0 1249.535 0.070 1249.605 ;
    RECT 0 1249.675 0.070 1249.745 ;
    RECT 0 1249.815 0.070 1249.885 ;
    RECT 0 1249.955 0.070 1250.025 ;
    RECT 0 1250.095 0.070 1250.165 ;
    RECT 0 1250.235 0.070 1250.305 ;
    RECT 0 1250.375 0.070 1250.445 ;
    RECT 0 1250.515 0.070 1250.585 ;
    RECT 0 1250.655 0.070 1250.725 ;
    RECT 0 1250.795 0.070 1250.865 ;
    RECT 0 1250.935 0.070 1251.005 ;
    RECT 0 1251.075 0.070 1251.145 ;
    RECT 0 1251.215 0.070 1251.285 ;
    RECT 0 1251.355 0.070 1251.425 ;
    RECT 0 1251.495 0.070 1251.565 ;
    RECT 0 1251.635 0.070 1251.705 ;
    RECT 0 1251.775 0.070 1251.845 ;
    RECT 0 1251.915 0.070 1251.985 ;
    RECT 0 1252.055 0.070 1252.125 ;
    RECT 0 1252.195 0.070 1252.265 ;
    RECT 0 1252.335 0.070 1252.405 ;
    RECT 0 1252.475 0.070 1252.545 ;
    RECT 0 1252.615 0.070 1252.685 ;
    RECT 0 1252.755 0.070 1252.825 ;
    RECT 0 1252.895 0.070 1252.965 ;
    RECT 0 1253.035 0.070 1253.105 ;
    RECT 0 1253.175 0.070 1253.245 ;
    RECT 0 1253.315 0.070 1253.385 ;
    RECT 0 1253.455 0.070 1253.525 ;
    RECT 0 1253.595 0.070 1253.665 ;
    RECT 0 1253.735 0.070 1253.805 ;
    RECT 0 1253.875 0.070 1253.945 ;
    RECT 0 1254.015 0.070 1254.085 ;
    RECT 0 1254.155 0.070 1254.225 ;
    RECT 0 1254.295 0.070 1254.365 ;
    RECT 0 1254.435 0.070 1254.505 ;
    RECT 0 1254.575 0.070 1254.645 ;
    RECT 0 1254.715 0.070 1254.785 ;
    RECT 0 1254.855 0.070 1254.925 ;
    RECT 0 1254.995 0.070 1255.065 ;
    RECT 0 1255.135 0.070 1255.205 ;
    RECT 0 1255.275 0.070 1255.345 ;
    RECT 0 1255.415 0.070 1255.485 ;
    RECT 0 1255.555 0.070 1255.625 ;
    RECT 0 1255.695 0.070 1255.765 ;
    RECT 0 1255.835 0.070 1255.905 ;
    RECT 0 1255.975 0.070 1256.045 ;
    RECT 0 1256.115 0.070 1256.185 ;
    RECT 0 1256.255 0.070 1256.325 ;
    RECT 0 1256.395 0.070 1256.465 ;
    RECT 0 1256.535 0.070 1256.605 ;
    RECT 0 1256.675 0.070 1256.745 ;
    RECT 0 1256.815 0.070 1256.885 ;
    RECT 0 1256.955 0.070 1257.025 ;
    RECT 0 1257.095 0.070 1257.165 ;
    RECT 0 1257.235 0.070 1257.305 ;
    RECT 0 1257.375 0.070 1257.445 ;
    RECT 0 1257.515 0.070 1257.585 ;
    RECT 0 1257.655 0.070 1257.725 ;
    RECT 0 1257.795 0.070 1257.865 ;
    RECT 0 1257.935 0.070 1258.005 ;
    RECT 0 1258.075 0.070 1258.145 ;
    RECT 0 1258.215 0.070 1258.285 ;
    RECT 0 1258.355 0.070 1258.425 ;
    RECT 0 1258.495 0.070 1258.565 ;
    RECT 0 1258.635 0.070 1258.705 ;
    RECT 0 1258.775 0.070 1258.845 ;
    RECT 0 1258.915 0.070 1258.985 ;
    RECT 0 1259.055 0.070 1259.125 ;
    RECT 0 1259.195 0.070 1259.265 ;
    RECT 0 1259.335 0.070 1259.405 ;
    RECT 0 1259.475 0.070 1259.545 ;
    RECT 0 1259.615 0.070 1259.685 ;
    RECT 0 1259.755 0.070 1259.825 ;
    RECT 0 1259.895 0.070 1259.965 ;
    RECT 0 1260.035 0.070 1260.105 ;
    RECT 0 1260.175 0.070 1260.245 ;
    RECT 0 1260.315 0.070 1260.385 ;
    RECT 0 1260.455 0.070 1260.525 ;
    RECT 0 1260.595 0.070 1260.665 ;
    RECT 0 1260.735 0.070 1260.805 ;
    RECT 0 1260.875 0.070 1260.945 ;
    RECT 0 1261.015 0.070 1261.085 ;
    RECT 0 1261.155 0.070 1261.225 ;
    RECT 0 1261.295 0.070 1261.365 ;
    RECT 0 1261.435 0.070 1261.505 ;
    RECT 0 1261.575 0.070 1261.645 ;
    RECT 0 1261.715 0.070 1261.785 ;
    RECT 0 1261.855 0.070 1261.925 ;
    RECT 0 1261.995 0.070 1262.065 ;
    RECT 0 1262.135 0.070 1262.205 ;
    RECT 0 1262.275 0.070 1262.345 ;
    RECT 0 1262.415 0.070 1262.485 ;
    RECT 0 1262.555 0.070 1262.625 ;
    RECT 0 1262.695 0.070 1262.765 ;
    RECT 0 1262.835 0.070 1262.905 ;
    RECT 0 1262.975 0.070 1263.045 ;
    RECT 0 1263.115 0.070 1263.185 ;
    RECT 0 1263.255 0.070 1263.325 ;
    RECT 0 1263.395 0.070 1263.465 ;
    RECT 0 1263.535 0.070 1263.605 ;
    RECT 0 1263.675 0.070 1263.745 ;
    RECT 0 1263.815 0.070 1263.885 ;
    RECT 0 1263.955 0.070 1264.025 ;
    RECT 0 1264.095 0.070 1264.165 ;
    RECT 0 1264.235 0.070 1264.305 ;
    RECT 0 1264.375 0.070 1264.445 ;
    RECT 0 1264.515 0.070 1264.585 ;
    RECT 0 1264.655 0.070 1264.725 ;
    RECT 0 1264.795 0.070 1264.865 ;
    RECT 0 1264.935 0.070 1265.005 ;
    RECT 0 1265.075 0.070 1265.145 ;
    RECT 0 1265.215 0.070 1265.285 ;
    RECT 0 1265.355 0.070 1265.425 ;
    RECT 0 1265.495 0.070 1265.565 ;
    RECT 0 1265.635 0.070 1265.705 ;
    RECT 0 1265.775 0.070 1265.845 ;
    RECT 0 1265.915 0.070 1265.985 ;
    RECT 0 1266.055 0.070 1266.125 ;
    RECT 0 1266.195 0.070 1266.265 ;
    RECT 0 1266.335 0.070 1266.405 ;
    RECT 0 1266.475 0.070 1266.545 ;
    RECT 0 1266.615 0.070 1266.685 ;
    RECT 0 1266.755 0.070 1266.825 ;
    RECT 0 1266.895 0.070 1266.965 ;
    RECT 0 1267.035 0.070 1267.105 ;
    RECT 0 1267.175 0.070 1267.245 ;
    RECT 0 1267.315 0.070 1267.385 ;
    RECT 0 1267.455 0.070 1267.525 ;
    RECT 0 1267.595 0.070 1267.665 ;
    RECT 0 1267.735 0.070 1267.805 ;
    RECT 0 1267.875 0.070 1267.945 ;
    RECT 0 1268.015 0.070 1268.085 ;
    RECT 0 1268.155 0.070 1268.225 ;
    RECT 0 1268.295 0.070 1268.365 ;
    RECT 0 1268.435 0.070 1268.505 ;
    RECT 0 1268.575 0.070 1268.645 ;
    RECT 0 1268.715 0.070 1268.785 ;
    RECT 0 1268.855 0.070 1268.925 ;
    RECT 0 1268.995 0.070 1269.065 ;
    RECT 0 1269.135 0.070 1269.205 ;
    RECT 0 1269.275 0.070 1269.345 ;
    RECT 0 1269.415 0.070 1269.485 ;
    RECT 0 1269.555 0.070 1269.625 ;
    RECT 0 1269.695 0.070 1269.765 ;
    RECT 0 1269.835 0.070 1269.905 ;
    RECT 0 1269.975 0.070 1270.045 ;
    RECT 0 1270.115 0.070 1270.185 ;
    RECT 0 1270.255 0.070 1270.325 ;
    RECT 0 1270.395 0.070 1270.465 ;
    RECT 0 1270.535 0.070 1270.605 ;
    RECT 0 1270.675 0.070 1270.745 ;
    RECT 0 1270.815 0.070 1270.885 ;
    RECT 0 1270.955 0.070 1271.025 ;
    RECT 0 1271.095 0.070 1271.165 ;
    RECT 0 1271.235 0.070 1271.305 ;
    RECT 0 1271.375 0.070 1271.445 ;
    RECT 0 1271.515 0.070 1271.585 ;
    RECT 0 1271.655 0.070 1271.725 ;
    RECT 0 1271.795 0.070 1271.865 ;
    RECT 0 1271.935 0.070 1272.005 ;
    RECT 0 1272.075 0.070 1272.145 ;
    RECT 0 1272.215 0.070 1272.285 ;
    RECT 0 1272.355 0.070 1272.425 ;
    RECT 0 1272.495 0.070 1272.565 ;
    RECT 0 1272.635 0.070 1272.705 ;
    RECT 0 1272.775 0.070 1272.845 ;
    RECT 0 1272.915 0.070 1272.985 ;
    RECT 0 1273.055 0.070 1273.125 ;
    RECT 0 1273.195 0.070 1273.265 ;
    RECT 0 1273.335 0.070 1273.405 ;
    RECT 0 1273.475 0.070 1273.545 ;
    RECT 0 1273.615 0.070 1273.685 ;
    RECT 0 1273.755 0.070 1273.825 ;
    RECT 0 1273.895 0.070 1273.965 ;
    RECT 0 1274.035 0.070 1274.105 ;
    RECT 0 1274.175 0.070 1274.245 ;
    RECT 0 1274.315 0.070 1274.385 ;
    RECT 0 1274.455 0.070 1274.525 ;
    RECT 0 1274.595 0.070 1274.665 ;
    RECT 0 1274.735 0.070 1274.805 ;
    RECT 0 1274.875 0.070 1274.945 ;
    RECT 0 1275.015 0.070 1275.085 ;
    RECT 0 1275.155 0.070 1275.225 ;
    RECT 0 1275.295 0.070 1275.365 ;
    RECT 0 1275.435 0.070 1275.505 ;
    RECT 0 1275.575 0.070 1275.645 ;
    RECT 0 1275.715 0.070 1275.785 ;
    RECT 0 1275.855 0.070 1275.925 ;
    RECT 0 1275.995 0.070 1276.065 ;
    RECT 0 1276.135 0.070 1276.205 ;
    RECT 0 1276.275 0.070 1276.345 ;
    RECT 0 1276.415 0.070 1276.485 ;
    RECT 0 1276.555 0.070 1276.625 ;
    RECT 0 1276.695 0.070 1276.765 ;
    RECT 0 1276.835 0.070 1276.905 ;
    RECT 0 1276.975 0.070 1277.045 ;
    RECT 0 1277.115 0.070 1277.185 ;
    RECT 0 1277.255 0.070 1277.325 ;
    RECT 0 1277.395 0.070 1277.465 ;
    RECT 0 1277.535 0.070 1277.605 ;
    RECT 0 1277.675 0.070 1277.745 ;
    RECT 0 1277.815 0.070 1277.885 ;
    RECT 0 1277.955 0.070 1278.025 ;
    RECT 0 1278.095 0.070 1278.165 ;
    RECT 0 1278.235 0.070 1278.305 ;
    RECT 0 1278.375 0.070 1278.445 ;
    RECT 0 1278.515 0.070 1278.585 ;
    RECT 0 1278.655 0.070 1278.725 ;
    RECT 0 1278.795 0.070 1278.865 ;
    RECT 0 1278.935 0.070 1279.005 ;
    RECT 0 1279.075 0.070 1279.145 ;
    RECT 0 1279.215 0.070 1279.285 ;
    RECT 0 1279.355 0.070 1279.425 ;
    RECT 0 1279.495 0.070 1279.565 ;
    RECT 0 1279.635 0.070 1279.705 ;
    RECT 0 1279.775 0.070 1279.845 ;
    RECT 0 1279.915 0.070 1279.985 ;
    RECT 0 1280.055 0.070 1280.125 ;
    RECT 0 1280.195 0.070 1280.265 ;
    RECT 0 1280.335 0.070 1280.405 ;
    RECT 0 1280.475 0.070 1280.545 ;
    RECT 0 1280.615 0.070 1280.685 ;
    RECT 0 1280.755 0.070 1280.825 ;
    RECT 0 1280.895 0.070 1280.965 ;
    RECT 0 1281.035 0.070 1281.105 ;
    RECT 0 1281.175 0.070 1281.245 ;
    RECT 0 1281.315 0.070 1281.385 ;
    RECT 0 1281.455 0.070 1281.525 ;
    RECT 0 1281.595 0.070 1281.665 ;
    RECT 0 1281.735 0.070 1281.805 ;
    RECT 0 1281.875 0.070 1281.945 ;
    RECT 0 1282.015 0.070 1282.085 ;
    RECT 0 1282.155 0.070 1282.225 ;
    RECT 0 1282.295 0.070 1282.365 ;
    RECT 0 1282.435 0.070 1282.505 ;
    RECT 0 1282.575 0.070 1282.645 ;
    RECT 0 1282.715 0.070 1282.785 ;
    RECT 0 1282.855 0.070 1282.925 ;
    RECT 0 1282.995 0.070 1283.065 ;
    RECT 0 1283.135 0.070 1283.205 ;
    RECT 0 1283.275 0.070 1283.345 ;
    RECT 0 1283.415 0.070 1283.485 ;
    RECT 0 1283.555 0.070 1283.625 ;
    RECT 0 1283.695 0.070 1283.765 ;
    RECT 0 1283.835 0.070 1283.905 ;
    RECT 0 1283.975 0.070 1284.045 ;
    RECT 0 1284.115 0.070 1284.185 ;
    RECT 0 1284.255 0.070 1284.325 ;
    RECT 0 1284.395 0.070 1284.465 ;
    RECT 0 1284.535 0.070 1284.605 ;
    RECT 0 1284.675 0.070 1284.745 ;
    RECT 0 1284.815 0.070 1284.885 ;
    RECT 0 1284.955 0.070 1285.025 ;
    RECT 0 1285.095 0.070 1285.165 ;
    RECT 0 1285.235 0.070 1285.305 ;
    RECT 0 1285.375 0.070 1285.445 ;
    RECT 0 1285.515 0.070 1285.585 ;
    RECT 0 1285.655 0.070 1285.725 ;
    RECT 0 1285.795 0.070 1285.865 ;
    RECT 0 1285.935 0.070 1286.005 ;
    RECT 0 1286.075 0.070 1286.145 ;
    RECT 0 1286.215 0.070 1286.285 ;
    RECT 0 1286.355 0.070 1286.425 ;
    RECT 0 1286.495 0.070 1286.565 ;
    RECT 0 1286.635 0.070 1286.705 ;
    RECT 0 1286.775 0.070 1286.845 ;
    RECT 0 1286.915 0.070 1286.985 ;
    RECT 0 1287.055 0.070 1287.125 ;
    RECT 0 1287.195 0.070 1287.265 ;
    RECT 0 1287.335 0.070 1287.405 ;
    RECT 0 1287.475 0.070 1287.545 ;
    RECT 0 1287.615 0.070 1287.685 ;
    RECT 0 1287.755 0.070 1287.825 ;
    RECT 0 1287.895 0.070 1287.965 ;
    RECT 0 1288.035 0.070 1288.105 ;
    RECT 0 1288.175 0.070 1288.245 ;
    RECT 0 1288.315 0.070 1288.385 ;
    RECT 0 1288.455 0.070 1288.525 ;
    RECT 0 1288.595 0.070 1288.665 ;
    RECT 0 1288.735 0.070 1288.805 ;
    RECT 0 1288.875 0.070 1288.945 ;
    RECT 0 1289.015 0.070 1289.085 ;
    RECT 0 1289.155 0.070 1289.225 ;
    RECT 0 1289.295 0.070 1289.365 ;
    RECT 0 1289.435 0.070 1289.505 ;
    RECT 0 1289.575 0.070 1289.645 ;
    RECT 0 1289.715 0.070 1289.785 ;
    RECT 0 1289.855 0.070 1289.925 ;
    RECT 0 1289.995 0.070 1290.065 ;
    RECT 0 1290.135 0.070 1290.205 ;
    RECT 0 1290.275 0.070 1290.345 ;
    RECT 0 1290.415 0.070 1290.485 ;
    RECT 0 1290.555 0.070 1290.625 ;
    RECT 0 1290.695 0.070 1290.765 ;
    RECT 0 1290.835 0.070 1290.905 ;
    RECT 0 1290.975 0.070 1291.045 ;
    RECT 0 1291.115 0.070 1291.185 ;
    RECT 0 1291.255 0.070 1291.325 ;
    RECT 0 1291.395 0.070 1291.465 ;
    RECT 0 1291.535 0.070 1291.605 ;
    RECT 0 1291.675 0.070 1291.745 ;
    RECT 0 1291.815 0.070 1291.885 ;
    RECT 0 1291.955 0.070 1292.025 ;
    RECT 0 1292.095 0.070 1292.165 ;
    RECT 0 1292.235 0.070 1292.305 ;
    RECT 0 1292.375 0.070 1292.445 ;
    RECT 0 1292.515 0.070 1292.585 ;
    RECT 0 1292.655 0.070 1292.725 ;
    RECT 0 1292.795 0.070 1292.865 ;
    RECT 0 1292.935 0.070 1293.005 ;
    RECT 0 1293.075 0.070 1293.145 ;
    RECT 0 1293.215 0.070 1293.285 ;
    RECT 0 1293.355 0.070 1293.425 ;
    RECT 0 1293.495 0.070 1293.565 ;
    RECT 0 1293.635 0.070 1293.705 ;
    RECT 0 1293.775 0.070 1293.845 ;
    RECT 0 1293.915 0.070 1293.985 ;
    RECT 0 1294.055 0.070 1294.125 ;
    RECT 0 1294.195 0.070 1294.265 ;
    RECT 0 1294.335 0.070 1294.405 ;
    RECT 0 1294.475 0.070 1294.545 ;
    RECT 0 1294.615 0.070 1294.685 ;
    RECT 0 1294.755 0.070 1294.825 ;
    RECT 0 1294.895 0.070 1294.965 ;
    RECT 0 1295.035 0.070 1295.105 ;
    RECT 0 1295.175 0.070 1295.245 ;
    RECT 0 1295.315 0.070 1295.385 ;
    RECT 0 1295.455 0.070 1295.525 ;
    RECT 0 1295.595 0.070 1295.665 ;
    RECT 0 1295.735 0.070 1295.805 ;
    RECT 0 1295.875 0.070 1295.945 ;
    RECT 0 1296.015 0.070 1296.085 ;
    RECT 0 1296.155 0.070 1296.225 ;
    RECT 0 1296.295 0.070 1296.365 ;
    RECT 0 1296.435 0.070 1296.505 ;
    RECT 0 1296.575 0.070 1296.645 ;
    RECT 0 1296.715 0.070 1296.785 ;
    RECT 0 1296.855 0.070 1296.925 ;
    RECT 0 1296.995 0.070 1297.065 ;
    RECT 0 1297.135 0.070 1297.205 ;
    RECT 0 1297.275 0.070 1297.345 ;
    RECT 0 1297.415 0.070 1297.485 ;
    RECT 0 1297.555 0.070 1297.625 ;
    RECT 0 1297.695 0.070 1297.765 ;
    RECT 0 1297.835 0.070 1297.905 ;
    RECT 0 1297.975 0.070 1298.045 ;
    RECT 0 1298.115 0.070 1298.185 ;
    RECT 0 1298.255 0.070 1298.325 ;
    RECT 0 1298.395 0.070 1298.465 ;
    RECT 0 1298.535 0.070 1298.605 ;
    RECT 0 1298.675 0.070 1298.745 ;
    RECT 0 1298.815 0.070 1298.885 ;
    RECT 0 1298.955 0.070 1299.025 ;
    RECT 0 1299.095 0.070 1299.165 ;
    RECT 0 1299.235 0.070 1299.305 ;
    RECT 0 1299.375 0.070 1299.445 ;
    RECT 0 1299.515 0.070 1299.585 ;
    RECT 0 1299.655 0.070 1299.725 ;
    RECT 0 1299.795 0.070 1299.865 ;
    RECT 0 1299.935 0.070 1300.005 ;
    RECT 0 1300.075 0.070 1300.145 ;
    RECT 0 1300.215 0.070 1300.285 ;
    RECT 0 1300.355 0.070 1300.425 ;
    RECT 0 1300.495 0.070 1300.565 ;
    RECT 0 1300.635 0.070 1300.705 ;
    RECT 0 1300.775 0.070 1300.845 ;
    RECT 0 1300.915 0.070 1300.985 ;
    RECT 0 1301.055 0.070 1301.125 ;
    RECT 0 1301.195 0.070 1301.265 ;
    RECT 0 1301.335 0.070 1301.405 ;
    RECT 0 1301.475 0.070 1301.545 ;
    RECT 0 1301.615 0.070 1301.685 ;
    RECT 0 1301.755 0.070 1301.825 ;
    RECT 0 1301.895 0.070 1301.965 ;
    RECT 0 1302.035 0.070 1302.105 ;
    RECT 0 1302.175 0.070 1302.245 ;
    RECT 0 1302.315 0.070 1302.385 ;
    RECT 0 1302.455 0.070 1302.525 ;
    RECT 0 1302.595 0.070 1302.665 ;
    RECT 0 1302.735 0.070 1302.805 ;
    RECT 0 1302.875 0.070 1302.945 ;
    RECT 0 1303.015 0.070 1303.085 ;
    RECT 0 1303.155 0.070 1303.225 ;
    RECT 0 1303.295 0.070 1303.365 ;
    RECT 0 1303.435 0.070 1303.505 ;
    RECT 0 1303.575 0.070 1303.645 ;
    RECT 0 1303.715 0.070 1303.785 ;
    RECT 0 1303.855 0.070 1303.925 ;
    RECT 0 1303.995 0.070 1304.065 ;
    RECT 0 1304.135 0.070 1304.205 ;
    RECT 0 1304.275 0.070 1304.345 ;
    RECT 0 1304.415 0.070 1304.485 ;
    RECT 0 1304.555 0.070 1304.625 ;
    RECT 0 1304.695 0.070 1304.765 ;
    RECT 0 1304.835 0.070 1304.905 ;
    RECT 0 1304.975 0.070 1305.045 ;
    RECT 0 1305.115 0.070 1305.185 ;
    RECT 0 1305.255 0.070 1305.325 ;
    RECT 0 1305.395 0.070 1305.465 ;
    RECT 0 1305.535 0.070 1305.605 ;
    RECT 0 1305.675 0.070 1305.745 ;
    RECT 0 1305.815 0.070 1305.885 ;
    RECT 0 1305.955 0.070 1306.025 ;
    RECT 0 1306.095 0.070 1306.165 ;
    RECT 0 1306.235 0.070 1306.305 ;
    RECT 0 1306.375 0.070 1306.445 ;
    RECT 0 1306.515 0.070 1306.585 ;
    RECT 0 1306.655 0.070 1306.725 ;
    RECT 0 1306.795 0.070 1306.865 ;
    RECT 0 1306.935 0.070 1307.005 ;
    RECT 0 1307.075 0.070 1307.145 ;
    RECT 0 1307.215 0.070 1307.285 ;
    RECT 0 1307.355 0.070 1307.425 ;
    RECT 0 1307.495 0.070 1307.565 ;
    RECT 0 1307.635 0.070 1307.705 ;
    RECT 0 1307.775 0.070 1307.845 ;
    RECT 0 1307.915 0.070 1307.985 ;
    RECT 0 1308.055 0.070 1308.125 ;
    RECT 0 1308.195 0.070 1308.265 ;
    RECT 0 1308.335 0.070 1308.405 ;
    RECT 0 1308.475 0.070 1308.545 ;
    RECT 0 1308.615 0.070 1308.685 ;
    RECT 0 1308.755 0.070 1308.825 ;
    RECT 0 1308.895 0.070 1308.965 ;
    RECT 0 1309.035 0.070 1309.105 ;
    RECT 0 1309.175 0.070 1309.245 ;
    RECT 0 1309.315 0.070 1309.385 ;
    RECT 0 1309.455 0.070 1309.525 ;
    RECT 0 1309.595 0.070 1309.665 ;
    RECT 0 1309.735 0.070 1309.805 ;
    RECT 0 1309.875 0.070 1309.945 ;
    RECT 0 1310.015 0.070 1310.085 ;
    RECT 0 1310.155 0.070 1310.225 ;
    RECT 0 1310.295 0.070 1310.365 ;
    RECT 0 1310.435 0.070 1310.505 ;
    RECT 0 1310.575 0.070 1310.645 ;
    RECT 0 1310.715 0.070 1310.785 ;
    RECT 0 1310.855 0.070 1310.925 ;
    RECT 0 1310.995 0.070 1311.065 ;
    RECT 0 1311.135 0.070 1311.205 ;
    RECT 0 1311.275 0.070 1311.345 ;
    RECT 0 1311.415 0.070 1311.485 ;
    RECT 0 1311.555 0.070 1311.625 ;
    RECT 0 1311.695 0.070 1311.765 ;
    RECT 0 1311.835 0.070 1311.905 ;
    RECT 0 1311.975 0.070 1312.045 ;
    RECT 0 1312.115 0.070 1312.185 ;
    RECT 0 1312.255 0.070 1312.325 ;
    RECT 0 1312.395 0.070 1312.465 ;
    RECT 0 1312.535 0.070 1312.605 ;
    RECT 0 1312.675 0.070 1312.745 ;
    RECT 0 1312.815 0.070 1312.885 ;
    RECT 0 1312.955 0.070 1313.025 ;
    RECT 0 1313.095 0.070 1313.165 ;
    RECT 0 1313.235 0.070 1313.305 ;
    RECT 0 1313.375 0.070 1313.445 ;
    RECT 0 1313.515 0.070 1313.585 ;
    RECT 0 1313.655 0.070 1313.725 ;
    RECT 0 1313.795 0.070 1313.865 ;
    RECT 0 1313.935 0.070 1314.005 ;
    RECT 0 1314.075 0.070 1314.145 ;
    RECT 0 1314.215 0.070 1314.285 ;
    RECT 0 1314.355 0.070 1314.425 ;
    RECT 0 1314.495 0.070 1314.565 ;
    RECT 0 1314.635 0.070 1314.705 ;
    RECT 0 1314.775 0.070 1314.845 ;
    RECT 0 1314.915 0.070 1314.985 ;
    RECT 0 1315.055 0.070 1315.125 ;
    RECT 0 1315.195 0.070 1315.265 ;
    RECT 0 1315.335 0.070 1315.405 ;
    RECT 0 1315.475 0.070 1315.545 ;
    RECT 0 1315.615 0.070 1315.685 ;
    RECT 0 1315.755 0.070 1315.825 ;
    RECT 0 1315.895 0.070 1315.965 ;
    RECT 0 1316.035 0.070 1316.105 ;
    RECT 0 1316.175 0.070 1316.245 ;
    RECT 0 1316.315 0.070 1316.385 ;
    RECT 0 1316.455 0.070 1316.525 ;
    RECT 0 1316.595 0.070 1316.665 ;
    RECT 0 1316.735 0.070 1316.805 ;
    RECT 0 1316.875 0.070 1316.945 ;
    RECT 0 1317.015 0.070 1317.085 ;
    RECT 0 1317.155 0.070 1317.225 ;
    RECT 0 1317.295 0.070 1317.365 ;
    RECT 0 1317.435 0.070 1317.505 ;
    RECT 0 1317.575 0.070 1317.645 ;
    RECT 0 1317.715 0.070 1317.785 ;
    RECT 0 1317.855 0.070 1317.925 ;
    RECT 0 1317.995 0.070 1318.065 ;
    RECT 0 1318.135 0.070 1318.205 ;
    RECT 0 1318.275 0.070 1318.345 ;
    RECT 0 1318.415 0.070 1318.485 ;
    RECT 0 1318.555 0.070 1318.625 ;
    RECT 0 1318.695 0.070 1318.765 ;
    RECT 0 1318.835 0.070 1318.905 ;
    RECT 0 1318.975 0.070 1319.045 ;
    RECT 0 1319.115 0.070 1319.185 ;
    RECT 0 1319.255 0.070 1319.325 ;
    RECT 0 1319.395 0.070 1319.465 ;
    RECT 0 1319.535 0.070 1319.605 ;
    RECT 0 1319.675 0.070 1319.745 ;
    RECT 0 1319.815 0.070 1319.885 ;
    RECT 0 1319.955 0.070 1320.025 ;
    RECT 0 1320.095 0.070 1320.165 ;
    RECT 0 1320.235 0.070 1320.305 ;
    RECT 0 1320.375 0.070 1320.445 ;
    RECT 0 1320.515 0.070 1320.585 ;
    RECT 0 1320.655 0.070 1320.725 ;
    RECT 0 1320.795 0.070 1320.865 ;
    RECT 0 1320.935 0.070 1321.005 ;
    RECT 0 1321.075 0.070 1321.145 ;
    RECT 0 1321.215 0.070 1321.285 ;
    RECT 0 1321.355 0.070 1321.425 ;
    RECT 0 1321.495 0.070 1321.565 ;
    RECT 0 1321.635 0.070 1321.705 ;
    RECT 0 1321.775 0.070 1321.845 ;
    RECT 0 1321.915 0.070 1321.985 ;
    RECT 0 1322.055 0.070 1322.125 ;
    RECT 0 1322.195 0.070 1322.265 ;
    RECT 0 1322.335 0.070 1322.405 ;
    RECT 0 1322.475 0.070 1322.545 ;
    RECT 0 1322.615 0.070 1322.685 ;
    RECT 0 1322.755 0.070 1322.825 ;
    RECT 0 1322.895 0.070 1322.965 ;
    RECT 0 1323.035 0.070 1323.105 ;
    RECT 0 1323.175 0.070 1323.245 ;
    RECT 0 1323.315 0.070 1323.385 ;
    RECT 0 1323.455 0.070 1323.525 ;
    RECT 0 1323.595 0.070 1323.665 ;
    RECT 0 1323.735 0.070 1323.805 ;
    RECT 0 1323.875 0.070 1323.945 ;
    RECT 0 1324.015 0.070 1324.085 ;
    RECT 0 1324.155 0.070 1324.225 ;
    RECT 0 1324.295 0.070 1324.365 ;
    RECT 0 1324.435 0.070 1324.505 ;
    RECT 0 1324.575 0.070 1324.645 ;
    RECT 0 1324.715 0.070 1324.785 ;
    RECT 0 1324.855 0.070 1324.925 ;
    RECT 0 1324.995 0.070 1325.065 ;
    RECT 0 1325.135 0.070 1325.205 ;
    RECT 0 1325.275 0.070 1325.345 ;
    RECT 0 1325.415 0.070 1325.485 ;
    RECT 0 1325.555 0.070 1325.625 ;
    RECT 0 1325.695 0.070 1325.765 ;
    RECT 0 1325.835 0.070 1325.905 ;
    RECT 0 1325.975 0.070 1326.045 ;
    RECT 0 1326.115 0.070 1326.185 ;
    RECT 0 1326.255 0.070 1326.325 ;
    RECT 0 1326.395 0.070 1326.465 ;
    RECT 0 1326.535 0.070 1326.605 ;
    RECT 0 1326.675 0.070 1326.745 ;
    RECT 0 1326.815 0.070 1326.885 ;
    RECT 0 1326.955 0.070 1327.025 ;
    RECT 0 1327.095 0.070 1327.165 ;
    RECT 0 1327.235 0.070 1327.305 ;
    RECT 0 1327.375 0.070 1327.445 ;
    RECT 0 1327.515 0.070 1327.585 ;
    RECT 0 1327.655 0.070 1327.725 ;
    RECT 0 1327.795 0.070 1327.865 ;
    RECT 0 1327.935 0.070 1328.005 ;
    RECT 0 1328.075 0.070 1328.145 ;
    RECT 0 1328.215 0.070 1328.285 ;
    RECT 0 1328.355 0.070 1328.425 ;
    RECT 0 1328.495 0.070 1328.565 ;
    RECT 0 1328.635 0.070 1328.705 ;
    RECT 0 1328.775 0.070 1328.845 ;
    RECT 0 1328.915 0.070 1328.985 ;
    RECT 0 1329.055 0.070 1329.125 ;
    RECT 0 1329.195 0.070 1329.265 ;
    RECT 0 1329.335 0.070 1329.405 ;
    RECT 0 1329.475 0.070 1329.545 ;
    RECT 0 1329.615 0.070 1329.685 ;
    RECT 0 1329.755 0.070 1329.825 ;
    RECT 0 1329.895 0.070 1329.965 ;
    RECT 0 1330.035 0.070 1330.105 ;
    RECT 0 1330.175 0.070 1330.245 ;
    RECT 0 1330.315 0.070 1330.385 ;
    RECT 0 1330.455 0.070 1330.525 ;
    RECT 0 1330.595 0.070 1330.665 ;
    RECT 0 1330.735 0.070 1330.805 ;
    RECT 0 1330.875 0.070 1330.945 ;
    RECT 0 1331.015 0.070 1331.085 ;
    RECT 0 1331.155 0.070 1331.225 ;
    RECT 0 1331.295 0.070 1331.365 ;
    RECT 0 1331.435 0.070 1331.505 ;
    RECT 0 1331.575 0.070 1331.645 ;
    RECT 0 1331.715 0.070 1331.785 ;
    RECT 0 1331.855 0.070 1331.925 ;
    RECT 0 1331.995 0.070 1332.065 ;
    RECT 0 1332.135 0.070 1332.205 ;
    RECT 0 1332.275 0.070 1332.345 ;
    RECT 0 1332.415 0.070 1332.485 ;
    RECT 0 1332.555 0.070 1332.625 ;
    RECT 0 1332.695 0.070 1332.765 ;
    RECT 0 1332.835 0.070 1332.905 ;
    RECT 0 1332.975 0.070 1333.045 ;
    RECT 0 1333.115 0.070 1333.185 ;
    RECT 0 1333.255 0.070 1333.325 ;
    RECT 0 1333.395 0.070 1333.465 ;
    RECT 0 1333.535 0.070 1333.605 ;
    RECT 0 1333.675 0.070 1333.745 ;
    RECT 0 1333.815 0.070 1333.885 ;
    RECT 0 1333.955 0.070 1334.025 ;
    RECT 0 1334.095 0.070 1334.165 ;
    RECT 0 1334.235 0.070 1334.305 ;
    RECT 0 1334.375 0.070 1334.445 ;
    RECT 0 1334.515 0.070 1334.585 ;
    RECT 0 1334.655 0.070 1334.725 ;
    RECT 0 1334.795 0.070 1334.865 ;
    RECT 0 1334.935 0.070 1335.005 ;
    RECT 0 1335.075 0.070 1335.145 ;
    RECT 0 1335.215 0.070 1335.285 ;
    RECT 0 1335.355 0.070 1335.425 ;
    RECT 0 1335.495 0.070 1335.565 ;
    RECT 0 1335.635 0.070 1335.705 ;
    RECT 0 1335.775 0.070 1335.845 ;
    RECT 0 1335.915 0.070 1335.985 ;
    RECT 0 1336.055 0.070 1336.125 ;
    RECT 0 1336.195 0.070 1336.265 ;
    RECT 0 1336.335 0.070 1336.405 ;
    RECT 0 1336.475 0.070 1336.545 ;
    RECT 0 1336.615 0.070 1336.685 ;
    RECT 0 1336.755 0.070 1336.825 ;
    RECT 0 1336.895 0.070 1336.965 ;
    RECT 0 1337.035 0.070 1337.105 ;
    RECT 0 1337.175 0.070 1337.245 ;
    RECT 0 1337.315 0.070 1337.385 ;
    RECT 0 1337.455 0.070 1337.525 ;
    RECT 0 1337.595 0.070 1337.665 ;
    RECT 0 1337.735 0.070 1337.805 ;
    RECT 0 1337.875 0.070 1337.945 ;
    RECT 0 1338.015 0.070 1338.085 ;
    RECT 0 1338.155 0.070 1338.225 ;
    RECT 0 1338.295 0.070 1338.365 ;
    RECT 0 1338.435 0.070 1338.505 ;
    RECT 0 1338.575 0.070 1338.645 ;
    RECT 0 1338.715 0.070 1338.785 ;
    RECT 0 1338.855 0.070 1338.925 ;
    RECT 0 1338.995 0.070 1339.065 ;
    RECT 0 1339.135 0.070 1339.205 ;
    RECT 0 1339.275 0.070 1339.345 ;
    RECT 0 1339.415 0.070 1339.485 ;
    RECT 0 1339.555 0.070 1339.625 ;
    RECT 0 1339.695 0.070 1339.765 ;
    RECT 0 1339.835 0.070 1339.905 ;
    RECT 0 1339.975 0.070 1340.045 ;
    RECT 0 1340.115 0.070 1340.185 ;
    RECT 0 1340.255 0.070 1340.325 ;
    RECT 0 1340.395 0.070 1340.465 ;
    RECT 0 1340.535 0.070 1340.605 ;
    RECT 0 1340.675 0.070 1340.745 ;
    RECT 0 1340.815 0.070 1340.885 ;
    RECT 0 1340.955 0.070 1341.025 ;
    RECT 0 1341.095 0.070 1341.165 ;
    RECT 0 1341.235 0.070 1341.305 ;
    RECT 0 1341.375 0.070 1341.445 ;
    RECT 0 1341.515 0.070 1341.585 ;
    RECT 0 1341.655 0.070 1341.725 ;
    RECT 0 1341.795 0.070 1341.865 ;
    RECT 0 1341.935 0.070 1342.005 ;
    RECT 0 1342.075 0.070 1342.145 ;
    RECT 0 1342.215 0.070 1342.285 ;
    RECT 0 1342.355 0.070 1342.425 ;
    RECT 0 1342.495 0.070 1342.565 ;
    RECT 0 1342.635 0.070 1342.705 ;
    RECT 0 1342.775 0.070 1342.845 ;
    RECT 0 1342.915 0.070 1342.985 ;
    RECT 0 1343.055 0.070 1343.125 ;
    RECT 0 1343.195 0.070 1343.265 ;
    RECT 0 1343.335 0.070 1343.405 ;
    RECT 0 1343.475 0.070 1343.545 ;
    RECT 0 1343.615 0.070 1343.685 ;
    RECT 0 1343.755 0.070 1343.825 ;
    RECT 0 1343.895 0.070 1343.965 ;
    RECT 0 1344.035 0.070 1344.105 ;
    RECT 0 1344.175 0.070 1344.245 ;
    RECT 0 1344.315 0.070 1344.385 ;
    RECT 0 1344.455 0.070 1344.525 ;
    RECT 0 1344.595 0.070 1344.665 ;
    RECT 0 1344.735 0.070 1344.805 ;
    RECT 0 1344.875 0.070 1344.945 ;
    RECT 0 1345.015 0.070 1345.085 ;
    RECT 0 1345.155 0.070 1345.225 ;
    RECT 0 1345.295 0.070 1345.365 ;
    RECT 0 1345.435 0.070 1345.505 ;
    RECT 0 1345.575 0.070 1345.645 ;
    RECT 0 1345.715 0.070 1345.785 ;
    RECT 0 1345.855 0.070 1345.925 ;
    RECT 0 1345.995 0.070 1346.065 ;
    RECT 0 1346.135 0.070 1346.205 ;
    RECT 0 1346.275 0.070 1346.345 ;
    RECT 0 1346.415 0.070 1346.485 ;
    RECT 0 1346.555 0.070 1346.625 ;
    RECT 0 1346.695 0.070 1346.765 ;
    RECT 0 1346.835 0.070 1346.905 ;
    RECT 0 1346.975 0.070 1347.045 ;
    RECT 0 1347.115 0.070 1347.185 ;
    RECT 0 1347.255 0.070 1347.325 ;
    RECT 0 1347.395 0.070 1347.465 ;
    RECT 0 1347.535 0.070 1347.605 ;
    RECT 0 1347.675 0.070 1347.745 ;
    RECT 0 1347.815 0.070 1347.885 ;
    RECT 0 1347.955 0.070 1348.025 ;
    RECT 0 1348.095 0.070 1348.165 ;
    RECT 0 1348.235 0.070 1348.305 ;
    RECT 0 1348.375 0.070 1348.445 ;
    RECT 0 1348.515 0.070 1348.585 ;
    RECT 0 1348.655 0.070 1348.725 ;
    RECT 0 1348.795 0.070 1348.865 ;
    RECT 0 1348.935 0.070 1349.005 ;
    RECT 0 1349.075 0.070 1349.145 ;
    RECT 0 1349.215 0.070 1349.285 ;
    RECT 0 1349.355 0.070 1349.425 ;
    RECT 0 1349.495 0.070 1349.565 ;
    RECT 0 1349.635 0.070 1349.705 ;
    RECT 0 1349.775 0.070 1349.845 ;
    RECT 0 1349.915 0.070 1349.985 ;
    RECT 0 1350.055 0.070 1350.125 ;
    RECT 0 1350.195 0.070 1350.265 ;
    RECT 0 1350.335 0.070 1350.405 ;
    RECT 0 1350.475 0.070 1350.545 ;
    RECT 0 1350.615 0.070 1350.685 ;
    RECT 0 1350.755 0.070 1350.825 ;
    RECT 0 1350.895 0.070 1350.965 ;
    RECT 0 1351.035 0.070 1351.105 ;
    RECT 0 1351.175 0.070 1351.245 ;
    RECT 0 1351.315 0.070 1351.385 ;
    RECT 0 1351.455 0.070 1351.525 ;
    RECT 0 1351.595 0.070 1351.665 ;
    RECT 0 1351.735 0.070 1351.805 ;
    RECT 0 1351.875 0.070 1351.945 ;
    RECT 0 1352.015 0.070 1352.085 ;
    RECT 0 1352.155 0.070 1352.225 ;
    RECT 0 1352.295 0.070 1352.365 ;
    RECT 0 1352.435 0.070 1352.505 ;
    RECT 0 1352.575 0.070 1352.645 ;
    RECT 0 1352.715 0.070 1352.785 ;
    RECT 0 1352.855 0.070 1352.925 ;
    RECT 0 1352.995 0.070 1353.065 ;
    RECT 0 1353.135 0.070 1353.205 ;
    RECT 0 1353.275 0.070 1353.345 ;
    RECT 0 1353.415 0.070 1353.485 ;
    RECT 0 1353.555 0.070 1353.625 ;
    RECT 0 1353.695 0.070 1353.765 ;
    RECT 0 1353.835 0.070 1353.905 ;
    RECT 0 1353.975 0.070 1354.045 ;
    RECT 0 1354.115 0.070 1354.185 ;
    RECT 0 1354.255 0.070 1354.325 ;
    RECT 0 1354.395 0.070 1354.465 ;
    RECT 0 1354.535 0.070 1354.605 ;
    RECT 0 1354.675 0.070 1354.745 ;
    RECT 0 1354.815 0.070 1354.885 ;
    RECT 0 1354.955 0.070 1355.025 ;
    RECT 0 1355.095 0.070 1355.165 ;
    RECT 0 1355.235 0.070 1355.305 ;
    RECT 0 1355.375 0.070 1355.445 ;
    RECT 0 1355.515 0.070 1355.585 ;
    RECT 0 1355.655 0.070 1355.725 ;
    RECT 0 1355.795 0.070 1355.865 ;
    RECT 0 1355.935 0.070 1356.005 ;
    RECT 0 1356.075 0.070 1356.145 ;
    RECT 0 1356.215 0.070 1356.285 ;
    RECT 0 1356.355 0.070 1356.425 ;
    RECT 0 1356.495 0.070 1356.565 ;
    RECT 0 1356.635 0.070 1356.705 ;
    RECT 0 1356.775 0.070 1356.845 ;
    RECT 0 1356.915 0.070 1356.985 ;
    RECT 0 1357.055 0.070 1357.125 ;
    RECT 0 1357.195 0.070 1357.265 ;
    RECT 0 1357.335 0.070 1357.405 ;
    RECT 0 1357.475 0.070 1357.545 ;
    RECT 0 1357.615 0.070 1357.685 ;
    RECT 0 1357.755 0.070 1357.825 ;
    RECT 0 1357.895 0.070 1357.965 ;
    RECT 0 1358.035 0.070 1358.105 ;
    RECT 0 1358.175 0.070 1358.245 ;
    RECT 0 1358.315 0.070 1358.385 ;
    RECT 0 1358.455 0.070 1358.525 ;
    RECT 0 1358.595 0.070 1358.665 ;
    RECT 0 1358.735 0.070 1358.805 ;
    RECT 0 1358.875 0.070 1358.945 ;
    RECT 0 1359.015 0.070 1359.085 ;
    RECT 0 1359.155 0.070 1359.225 ;
    RECT 0 1359.295 0.070 1359.365 ;
    RECT 0 1359.435 0.070 1359.505 ;
    RECT 0 1359.575 0.070 1359.645 ;
    RECT 0 1359.715 0.070 1359.785 ;
    RECT 0 1359.855 0.070 1359.925 ;
    RECT 0 1359.995 0.070 1360.065 ;
    RECT 0 1360.135 0.070 1360.205 ;
    RECT 0 1360.275 0.070 1360.345 ;
    RECT 0 1360.415 0.070 1360.485 ;
    RECT 0 1360.555 0.070 1360.625 ;
    RECT 0 1360.695 0.070 1360.765 ;
    RECT 0 1360.835 0.070 1360.905 ;
    RECT 0 1360.975 0.070 1361.045 ;
    RECT 0 1361.115 0.070 1361.185 ;
    RECT 0 1361.255 0.070 1361.325 ;
    RECT 0 1361.395 0.070 1361.465 ;
    RECT 0 1361.535 0.070 1361.605 ;
    RECT 0 1361.675 0.070 1361.745 ;
    RECT 0 1361.815 0.070 1361.885 ;
    RECT 0 1361.955 0.070 1362.025 ;
    RECT 0 1362.095 0.070 1362.165 ;
    RECT 0 1362.235 0.070 1362.305 ;
    RECT 0 1362.375 0.070 1362.445 ;
    RECT 0 1362.515 0.070 1362.585 ;
    RECT 0 1362.655 0.070 1362.725 ;
    RECT 0 1362.795 0.070 1362.865 ;
    RECT 0 1362.935 0.070 1363.005 ;
    RECT 0 1363.075 0.070 1363.145 ;
    RECT 0 1363.215 0.070 1363.285 ;
    RECT 0 1363.355 0.070 1363.425 ;
    RECT 0 1363.495 0.070 1363.565 ;
    RECT 0 1363.635 0.070 1363.705 ;
    RECT 0 1363.775 0.070 1363.845 ;
    RECT 0 1363.915 0.070 1363.985 ;
    RECT 0 1364.055 0.070 1364.125 ;
    RECT 0 1364.195 0.070 1364.265 ;
    RECT 0 1364.335 0.070 1364.405 ;
    RECT 0 1364.475 0.070 1364.545 ;
    RECT 0 1364.615 0.070 1364.685 ;
    RECT 0 1364.755 0.070 1364.825 ;
    RECT 0 1364.895 0.070 1364.965 ;
    RECT 0 1365.035 0.070 1365.105 ;
    RECT 0 1365.175 0.070 1365.245 ;
    RECT 0 1365.315 0.070 1365.385 ;
    RECT 0 1365.455 0.070 1365.525 ;
    RECT 0 1365.595 0.070 1365.665 ;
    RECT 0 1365.735 0.070 1365.805 ;
    RECT 0 1365.875 0.070 1365.945 ;
    RECT 0 1366.015 0.070 1366.085 ;
    RECT 0 1366.155 0.070 1366.225 ;
    RECT 0 1366.295 0.070 1366.365 ;
    RECT 0 1366.435 0.070 1366.505 ;
    RECT 0 1366.575 0.070 1366.645 ;
    RECT 0 1366.715 0.070 1366.785 ;
    RECT 0 1366.855 0.070 1366.925 ;
    RECT 0 1366.995 0.070 1367.065 ;
    RECT 0 1367.135 0.070 1367.205 ;
    RECT 0 1367.275 0.070 1367.345 ;
    RECT 0 1367.415 0.070 1367.485 ;
    RECT 0 1367.555 0.070 1367.625 ;
    RECT 0 1367.695 0.070 1367.765 ;
    RECT 0 1367.835 0.070 1367.905 ;
    RECT 0 1367.975 0.070 1368.045 ;
    RECT 0 1368.115 0.070 1368.185 ;
    RECT 0 1368.255 0.070 1368.325 ;
    RECT 0 1368.395 0.070 1368.465 ;
    RECT 0 1368.535 0.070 1368.605 ;
    RECT 0 1368.675 0.070 1368.745 ;
    RECT 0 1368.815 0.070 1368.885 ;
    RECT 0 1368.955 0.070 1369.025 ;
    RECT 0 1369.095 0.070 1369.165 ;
    RECT 0 1369.235 0.070 1369.305 ;
    RECT 0 1369.375 0.070 1369.445 ;
    RECT 0 1369.515 0.070 1369.585 ;
    RECT 0 1369.655 0.070 1369.725 ;
    RECT 0 1369.795 0.070 1369.865 ;
    RECT 0 1369.935 0.070 1370.005 ;
    RECT 0 1370.075 0.070 1370.145 ;
    RECT 0 1370.215 0.070 1370.285 ;
    RECT 0 1370.355 0.070 1370.425 ;
    RECT 0 1370.495 0.070 1370.565 ;
    RECT 0 1370.635 0.070 1370.705 ;
    RECT 0 1370.775 0.070 1370.845 ;
    RECT 0 1370.915 0.070 1370.985 ;
    RECT 0 1371.055 0.070 1371.125 ;
    RECT 0 1371.195 0.070 1371.265 ;
    RECT 0 1371.335 0.070 1371.405 ;
    RECT 0 1371.475 0.070 1371.545 ;
    RECT 0 1371.615 0.070 1371.685 ;
    RECT 0 1371.755 0.070 1371.825 ;
    RECT 0 1371.895 0.070 1371.965 ;
    RECT 0 1372.035 0.070 1372.105 ;
    RECT 0 1372.175 0.070 1372.245 ;
    RECT 0 1372.315 0.070 1372.385 ;
    RECT 0 1372.455 0.070 1372.525 ;
    RECT 0 1372.595 0.070 1372.665 ;
    RECT 0 1372.735 0.070 1372.805 ;
    RECT 0 1372.875 0.070 1372.945 ;
    RECT 0 1373.015 0.070 1373.085 ;
    RECT 0 1373.155 0.070 1373.225 ;
    RECT 0 1373.295 0.070 1373.365 ;
    RECT 0 1373.435 0.070 1373.505 ;
    RECT 0 1373.575 0.070 1373.645 ;
    RECT 0 1373.715 0.070 1373.785 ;
    RECT 0 1373.855 0.070 1373.925 ;
    RECT 0 1373.995 0.070 1374.065 ;
    RECT 0 1374.135 0.070 1374.205 ;
    RECT 0 1374.275 0.070 1374.345 ;
    RECT 0 1374.415 0.070 1374.485 ;
    RECT 0 1374.555 0.070 1374.625 ;
    RECT 0 1374.695 0.070 1374.765 ;
    RECT 0 1374.835 0.070 1374.905 ;
    RECT 0 1374.975 0.070 1375.045 ;
    RECT 0 1375.115 0.070 1375.185 ;
    RECT 0 1375.255 0.070 1375.325 ;
    RECT 0 1375.395 0.070 1375.465 ;
    RECT 0 1375.535 0.070 1375.605 ;
    RECT 0 1375.675 0.070 1375.745 ;
    RECT 0 1375.815 0.070 1375.885 ;
    RECT 0 1375.955 0.070 1376.025 ;
    RECT 0 1376.095 0.070 1376.165 ;
    RECT 0 1376.235 0.070 1376.305 ;
    RECT 0 1376.375 0.070 1376.445 ;
    RECT 0 1376.515 0.070 1376.585 ;
    RECT 0 1376.655 0.070 1376.725 ;
    RECT 0 1376.795 0.070 1376.865 ;
    RECT 0 1376.935 0.070 1377.005 ;
    RECT 0 1377.075 0.070 1377.145 ;
    RECT 0 1377.215 0.070 1377.285 ;
    RECT 0 1377.355 0.070 1377.425 ;
    RECT 0 1377.495 0.070 1377.565 ;
    RECT 0 1377.635 0.070 1377.705 ;
    RECT 0 1377.775 0.070 1377.845 ;
    RECT 0 1377.915 0.070 1377.985 ;
    RECT 0 1378.055 0.070 1378.125 ;
    RECT 0 1378.195 0.070 1378.265 ;
    RECT 0 1378.335 0.070 1378.405 ;
    RECT 0 1378.475 0.070 1378.545 ;
    RECT 0 1378.615 0.070 1378.685 ;
    RECT 0 1378.755 0.070 1378.825 ;
    RECT 0 1378.895 0.070 1378.965 ;
    RECT 0 1379.035 0.070 1379.105 ;
    RECT 0 1379.175 0.070 1379.245 ;
    RECT 0 1379.315 0.070 1379.385 ;
    RECT 0 1379.455 0.070 1379.525 ;
    RECT 0 1379.595 0.070 1379.665 ;
    RECT 0 1379.735 0.070 1379.805 ;
    RECT 0 1379.875 0.070 1379.945 ;
    RECT 0 1380.015 0.070 1380.085 ;
    RECT 0 1380.155 0.070 1380.225 ;
    RECT 0 1380.295 0.070 1380.365 ;
    RECT 0 1380.435 0.070 1380.505 ;
    RECT 0 1380.575 0.070 1380.645 ;
    RECT 0 1380.715 0.070 1380.785 ;
    RECT 0 1380.855 0.070 1380.925 ;
    RECT 0 1380.995 0.070 1381.065 ;
    RECT 0 1381.135 0.070 1381.205 ;
    RECT 0 1381.275 0.070 1381.345 ;
    RECT 0 1381.415 0.070 1381.485 ;
    RECT 0 1381.555 0.070 1381.625 ;
    RECT 0 1381.695 0.070 1381.765 ;
    RECT 0 1381.835 0.070 1381.905 ;
    RECT 0 1381.975 0.070 1382.045 ;
    RECT 0 1382.115 0.070 1382.185 ;
    RECT 0 1382.255 0.070 1382.325 ;
    RECT 0 1382.395 0.070 1382.465 ;
    RECT 0 1382.535 0.070 1382.605 ;
    RECT 0 1382.675 0.070 1382.745 ;
    RECT 0 1382.815 0.070 1382.885 ;
    RECT 0 1382.955 0.070 1383.025 ;
    RECT 0 1383.095 0.070 1383.165 ;
    RECT 0 1383.235 0.070 1383.305 ;
    RECT 0 1383.375 0.070 1383.445 ;
    RECT 0 1383.515 0.070 1383.585 ;
    RECT 0 1383.655 0.070 1383.725 ;
    RECT 0 1383.795 0.070 1383.865 ;
    RECT 0 1383.935 0.070 1384.005 ;
    RECT 0 1384.075 0.070 1384.145 ;
    RECT 0 1384.215 0.070 1384.285 ;
    RECT 0 1384.355 0.070 1384.425 ;
    RECT 0 1384.495 0.070 1384.565 ;
    RECT 0 1384.635 0.070 1384.705 ;
    RECT 0 1384.775 0.070 1384.845 ;
    RECT 0 1384.915 0.070 1384.985 ;
    RECT 0 1385.055 0.070 1385.125 ;
    RECT 0 1385.195 0.070 1385.265 ;
    RECT 0 1385.335 0.070 1385.405 ;
    RECT 0 1385.475 0.070 1385.545 ;
    RECT 0 1385.615 0.070 1385.685 ;
    RECT 0 1385.755 0.070 1385.825 ;
    RECT 0 1385.895 0.070 1385.965 ;
    RECT 0 1386.035 0.070 1386.105 ;
    RECT 0 1386.175 0.070 1386.245 ;
    RECT 0 1386.315 0.070 1386.385 ;
    RECT 0 1386.455 0.070 1386.525 ;
    RECT 0 1386.595 0.070 1386.665 ;
    RECT 0 1386.735 0.070 1386.805 ;
    RECT 0 1386.875 0.070 1386.945 ;
    RECT 0 1387.015 0.070 1387.085 ;
    RECT 0 1387.155 0.070 1387.225 ;
    RECT 0 1387.295 0.070 1387.365 ;
    RECT 0 1387.435 0.070 1387.505 ;
    RECT 0 1387.575 0.070 1387.645 ;
    RECT 0 1387.715 0.070 1387.785 ;
    RECT 0 1387.855 0.070 1387.925 ;
    RECT 0 1387.995 0.070 1388.065 ;
    RECT 0 1388.135 0.070 1388.205 ;
    RECT 0 1388.275 0.070 1388.345 ;
    RECT 0 1388.415 0.070 1388.485 ;
    RECT 0 1388.555 0.070 1388.625 ;
    RECT 0 1388.695 0.070 1388.765 ;
    RECT 0 1388.835 0.070 1388.905 ;
    RECT 0 1388.975 0.070 1389.045 ;
    RECT 0 1389.115 0.070 1389.185 ;
    RECT 0 1389.255 0.070 1389.325 ;
    RECT 0 1389.395 0.070 1389.465 ;
    RECT 0 1389.535 0.070 1389.605 ;
    RECT 0 1389.675 0.070 1389.745 ;
    RECT 0 1389.815 0.070 1389.885 ;
    RECT 0 1389.955 0.070 1390.025 ;
    RECT 0 1390.095 0.070 1390.165 ;
    RECT 0 1390.235 0.070 1390.305 ;
    RECT 0 1390.375 0.070 1390.445 ;
    RECT 0 1390.515 0.070 1390.585 ;
    RECT 0 1390.655 0.070 1390.725 ;
    RECT 0 1390.795 0.070 1390.865 ;
    RECT 0 1390.935 0.070 1391.005 ;
    RECT 0 1391.075 0.070 1391.145 ;
    RECT 0 1391.215 0.070 1391.285 ;
    RECT 0 1391.355 0.070 1391.425 ;
    RECT 0 1391.495 0.070 1391.565 ;
    RECT 0 1391.635 0.070 1391.705 ;
    RECT 0 1391.775 0.070 1391.845 ;
    RECT 0 1391.915 0.070 1391.985 ;
    RECT 0 1392.055 0.070 1392.125 ;
    RECT 0 1392.195 0.070 1392.265 ;
    RECT 0 1392.335 0.070 1392.405 ;
    RECT 0 1392.475 0.070 1392.545 ;
    RECT 0 1392.615 0.070 1392.685 ;
    RECT 0 1392.755 0.070 1392.825 ;
    RECT 0 1392.895 0.070 1392.965 ;
    RECT 0 1393.035 0.070 1393.105 ;
    RECT 0 1393.175 0.070 1393.245 ;
    RECT 0 1393.315 0.070 1393.385 ;
    RECT 0 1393.455 0.070 1393.525 ;
    RECT 0 1393.595 0.070 1393.665 ;
    RECT 0 1393.735 0.070 1393.805 ;
    RECT 0 1393.875 0.070 1393.945 ;
    RECT 0 1394.015 0.070 1394.085 ;
    RECT 0 1394.155 0.070 1394.225 ;
    RECT 0 1394.295 0.070 1394.365 ;
    RECT 0 1394.435 0.070 1394.505 ;
    RECT 0 1394.575 0.070 1394.645 ;
    RECT 0 1394.715 0.070 1394.785 ;
    RECT 0 1394.855 0.070 1394.925 ;
    RECT 0 1394.995 0.070 1395.065 ;
    RECT 0 1395.135 0.070 1395.205 ;
    RECT 0 1395.275 0.070 1395.345 ;
    RECT 0 1395.415 0.070 1395.485 ;
    RECT 0 1395.555 0.070 1395.625 ;
    RECT 0 1395.695 0.070 1395.765 ;
    RECT 0 1395.835 0.070 1395.905 ;
    RECT 0 1395.975 0.070 1396.045 ;
    RECT 0 1396.115 0.070 1396.185 ;
    RECT 0 1396.255 0.070 1396.325 ;
    RECT 0 1396.395 0.070 1396.465 ;
    RECT 0 1396.535 0.070 1396.605 ;
    RECT 0 1396.675 0.070 1396.745 ;
    RECT 0 1396.815 0.070 1396.885 ;
    RECT 0 1396.955 0.070 1397.025 ;
    RECT 0 1397.095 0.070 1397.165 ;
    RECT 0 1397.235 0.070 1397.305 ;
    RECT 0 1397.375 0.070 1397.445 ;
    RECT 0 1397.515 0.070 1397.585 ;
    RECT 0 1397.655 0.070 1397.725 ;
    RECT 0 1397.795 0.070 1397.865 ;
    RECT 0 1397.935 0.070 1398.005 ;
    RECT 0 1398.075 0.070 1398.145 ;
    RECT 0 1398.215 0.070 1398.285 ;
    RECT 0 1398.355 0.070 1398.425 ;
    RECT 0 1398.495 0.070 1398.565 ;
    RECT 0 1398.635 0.070 1398.705 ;
    RECT 0 1398.775 0.070 1398.845 ;
    RECT 0 1398.915 0.070 1398.985 ;
    RECT 0 1399.055 0.070 1399.125 ;
    RECT 0 1399.195 0.070 1399.265 ;
    RECT 0 1399.335 0.070 1399.405 ;
    RECT 0 1399.475 0.070 1399.545 ;
    RECT 0 1399.615 0.070 1399.685 ;
    RECT 0 1399.755 0.070 1399.825 ;
    RECT 0 1399.895 0.070 1399.965 ;
    RECT 0 1400.035 0.070 1400.105 ;
    RECT 0 1400.175 0.070 1400.245 ;
    RECT 0 1400.315 0.070 1400.385 ;
    RECT 0 1400.455 0.070 1400.525 ;
    RECT 0 1400.595 0.070 1400.665 ;
    RECT 0 1400.735 0.070 1400.805 ;
    RECT 0 1400.875 0.070 1400.945 ;
    RECT 0 1401.015 0.070 1401.085 ;
    RECT 0 1401.155 0.070 1401.225 ;
    RECT 0 1401.295 0.070 1401.365 ;
    RECT 0 1401.435 0.070 1401.505 ;
    RECT 0 1401.575 0.070 1401.645 ;
    RECT 0 1401.715 0.070 1401.785 ;
    RECT 0 1401.855 0.070 1401.925 ;
    RECT 0 1401.995 0.070 1402.065 ;
    RECT 0 1402.135 0.070 1402.205 ;
    RECT 0 1402.275 0.070 1402.345 ;
    RECT 0 1402.415 0.070 1402.485 ;
    RECT 0 1402.555 0.070 1402.625 ;
    RECT 0 1402.695 0.070 1402.765 ;
    RECT 0 1402.835 0.070 1402.905 ;
    RECT 0 1402.975 0.070 1403.045 ;
    RECT 0 1403.115 0.070 1403.185 ;
    RECT 0 1403.255 0.070 1403.325 ;
    RECT 0 1403.395 0.070 1403.465 ;
    RECT 0 1403.535 0.070 1403.605 ;
    RECT 0 1403.675 0.070 1403.745 ;
    RECT 0 1403.815 0.070 1403.885 ;
    RECT 0 1403.955 0.070 1404.025 ;
    RECT 0 1404.095 0.070 1404.165 ;
    RECT 0 1404.235 0.070 1404.305 ;
    RECT 0 1404.375 0.070 1404.445 ;
    RECT 0 1404.515 0.070 1404.585 ;
    RECT 0 1404.655 0.070 1404.725 ;
    RECT 0 1404.795 0.070 1404.865 ;
    RECT 0 1404.935 0.070 1405.005 ;
    RECT 0 1405.075 0.070 1405.145 ;
    RECT 0 1405.215 0.070 1405.285 ;
    RECT 0 1405.355 0.070 1405.425 ;
    RECT 0 1405.495 0.070 1405.565 ;
    RECT 0 1405.635 0.070 1405.705 ;
    RECT 0 1405.775 0.070 1405.845 ;
    RECT 0 1405.915 0.070 1405.985 ;
    RECT 0 1406.055 0.070 1406.125 ;
    RECT 0 1406.195 0.070 1406.265 ;
    RECT 0 1406.335 0.070 1510.845 ;
    RECT 0 1510.915 0.070 1510.985 ;
    RECT 0 1511.055 0.070 1511.125 ;
    RECT 0 1511.195 0.070 1511.265 ;
    RECT 0 1511.335 0.070 1511.405 ;
    RECT 0 1511.475 0.070 1615.985 ;
    RECT 0 1616.055 0.070 1616.125 ;
    RECT 0 1616.195 0.070 1616.265 ;
    RECT 0 1616.335 0.070 1618.400 ;
    LAYER metal4 ;
    RECT 0 0 2078.600 1.400 ;
    RECT 0 1617.000 2078.600 1618.400 ;
    RECT 0.000 1.400 1.260 1617.000 ;
    RECT 1.540 1.400 2.380 1617.000 ;
    RECT 2.660 1.400 3.500 1617.000 ;
    RECT 3.780 1.400 4.620 1617.000 ;
    RECT 4.900 1.400 5.740 1617.000 ;
    RECT 6.020 1.400 6.860 1617.000 ;
    RECT 7.140 1.400 7.980 1617.000 ;
    RECT 8.260 1.400 9.100 1617.000 ;
    RECT 9.380 1.400 10.220 1617.000 ;
    RECT 10.500 1.400 11.340 1617.000 ;
    RECT 11.620 1.400 12.460 1617.000 ;
    RECT 12.740 1.400 13.580 1617.000 ;
    RECT 13.860 1.400 14.700 1617.000 ;
    RECT 14.980 1.400 15.820 1617.000 ;
    RECT 16.100 1.400 16.940 1617.000 ;
    RECT 17.220 1.400 18.060 1617.000 ;
    RECT 18.340 1.400 19.180 1617.000 ;
    RECT 19.460 1.400 20.300 1617.000 ;
    RECT 20.580 1.400 21.420 1617.000 ;
    RECT 21.700 1.400 22.540 1617.000 ;
    RECT 22.820 1.400 23.660 1617.000 ;
    RECT 23.940 1.400 24.780 1617.000 ;
    RECT 25.060 1.400 25.900 1617.000 ;
    RECT 26.180 1.400 27.020 1617.000 ;
    RECT 27.300 1.400 28.140 1617.000 ;
    RECT 28.420 1.400 29.260 1617.000 ;
    RECT 29.540 1.400 30.380 1617.000 ;
    RECT 30.660 1.400 31.500 1617.000 ;
    RECT 31.780 1.400 32.620 1617.000 ;
    RECT 32.900 1.400 33.740 1617.000 ;
    RECT 34.020 1.400 34.860 1617.000 ;
    RECT 35.140 1.400 35.980 1617.000 ;
    RECT 36.260 1.400 37.100 1617.000 ;
    RECT 37.380 1.400 38.220 1617.000 ;
    RECT 38.500 1.400 39.340 1617.000 ;
    RECT 39.620 1.400 40.460 1617.000 ;
    RECT 40.740 1.400 41.580 1617.000 ;
    RECT 41.860 1.400 42.700 1617.000 ;
    RECT 42.980 1.400 43.820 1617.000 ;
    RECT 44.100 1.400 44.940 1617.000 ;
    RECT 45.220 1.400 46.060 1617.000 ;
    RECT 46.340 1.400 47.180 1617.000 ;
    RECT 47.460 1.400 48.300 1617.000 ;
    RECT 48.580 1.400 49.420 1617.000 ;
    RECT 49.700 1.400 50.540 1617.000 ;
    RECT 50.820 1.400 51.660 1617.000 ;
    RECT 51.940 1.400 52.780 1617.000 ;
    RECT 53.060 1.400 53.900 1617.000 ;
    RECT 54.180 1.400 55.020 1617.000 ;
    RECT 55.300 1.400 56.140 1617.000 ;
    RECT 56.420 1.400 57.260 1617.000 ;
    RECT 57.540 1.400 58.380 1617.000 ;
    RECT 58.660 1.400 59.500 1617.000 ;
    RECT 59.780 1.400 60.620 1617.000 ;
    RECT 60.900 1.400 61.740 1617.000 ;
    RECT 62.020 1.400 62.860 1617.000 ;
    RECT 63.140 1.400 63.980 1617.000 ;
    RECT 64.260 1.400 65.100 1617.000 ;
    RECT 65.380 1.400 66.220 1617.000 ;
    RECT 66.500 1.400 67.340 1617.000 ;
    RECT 67.620 1.400 68.460 1617.000 ;
    RECT 68.740 1.400 69.580 1617.000 ;
    RECT 69.860 1.400 70.700 1617.000 ;
    RECT 70.980 1.400 71.820 1617.000 ;
    RECT 72.100 1.400 72.940 1617.000 ;
    RECT 73.220 1.400 74.060 1617.000 ;
    RECT 74.340 1.400 75.180 1617.000 ;
    RECT 75.460 1.400 76.300 1617.000 ;
    RECT 76.580 1.400 77.420 1617.000 ;
    RECT 77.700 1.400 78.540 1617.000 ;
    RECT 78.820 1.400 79.660 1617.000 ;
    RECT 79.940 1.400 80.780 1617.000 ;
    RECT 81.060 1.400 81.900 1617.000 ;
    RECT 82.180 1.400 83.020 1617.000 ;
    RECT 83.300 1.400 84.140 1617.000 ;
    RECT 84.420 1.400 85.260 1617.000 ;
    RECT 85.540 1.400 86.380 1617.000 ;
    RECT 86.660 1.400 87.500 1617.000 ;
    RECT 87.780 1.400 88.620 1617.000 ;
    RECT 88.900 1.400 89.740 1617.000 ;
    RECT 90.020 1.400 90.860 1617.000 ;
    RECT 91.140 1.400 91.980 1617.000 ;
    RECT 92.260 1.400 93.100 1617.000 ;
    RECT 93.380 1.400 94.220 1617.000 ;
    RECT 94.500 1.400 95.340 1617.000 ;
    RECT 95.620 1.400 96.460 1617.000 ;
    RECT 96.740 1.400 97.580 1617.000 ;
    RECT 97.860 1.400 98.700 1617.000 ;
    RECT 98.980 1.400 99.820 1617.000 ;
    RECT 100.100 1.400 100.940 1617.000 ;
    RECT 101.220 1.400 102.060 1617.000 ;
    RECT 102.340 1.400 103.180 1617.000 ;
    RECT 103.460 1.400 104.300 1617.000 ;
    RECT 104.580 1.400 105.420 1617.000 ;
    RECT 105.700 1.400 106.540 1617.000 ;
    RECT 106.820 1.400 107.660 1617.000 ;
    RECT 107.940 1.400 108.780 1617.000 ;
    RECT 109.060 1.400 109.900 1617.000 ;
    RECT 110.180 1.400 111.020 1617.000 ;
    RECT 111.300 1.400 112.140 1617.000 ;
    RECT 112.420 1.400 113.260 1617.000 ;
    RECT 113.540 1.400 114.380 1617.000 ;
    RECT 114.660 1.400 115.500 1617.000 ;
    RECT 115.780 1.400 116.620 1617.000 ;
    RECT 116.900 1.400 117.740 1617.000 ;
    RECT 118.020 1.400 118.860 1617.000 ;
    RECT 119.140 1.400 119.980 1617.000 ;
    RECT 120.260 1.400 121.100 1617.000 ;
    RECT 121.380 1.400 122.220 1617.000 ;
    RECT 122.500 1.400 123.340 1617.000 ;
    RECT 123.620 1.400 124.460 1617.000 ;
    RECT 124.740 1.400 125.580 1617.000 ;
    RECT 125.860 1.400 126.700 1617.000 ;
    RECT 126.980 1.400 127.820 1617.000 ;
    RECT 128.100 1.400 128.940 1617.000 ;
    RECT 129.220 1.400 130.060 1617.000 ;
    RECT 130.340 1.400 131.180 1617.000 ;
    RECT 131.460 1.400 132.300 1617.000 ;
    RECT 132.580 1.400 133.420 1617.000 ;
    RECT 133.700 1.400 134.540 1617.000 ;
    RECT 134.820 1.400 135.660 1617.000 ;
    RECT 135.940 1.400 136.780 1617.000 ;
    RECT 137.060 1.400 137.900 1617.000 ;
    RECT 138.180 1.400 139.020 1617.000 ;
    RECT 139.300 1.400 140.140 1617.000 ;
    RECT 140.420 1.400 141.260 1617.000 ;
    RECT 141.540 1.400 142.380 1617.000 ;
    RECT 142.660 1.400 143.500 1617.000 ;
    RECT 143.780 1.400 144.620 1617.000 ;
    RECT 144.900 1.400 145.740 1617.000 ;
    RECT 146.020 1.400 146.860 1617.000 ;
    RECT 147.140 1.400 147.980 1617.000 ;
    RECT 148.260 1.400 149.100 1617.000 ;
    RECT 149.380 1.400 150.220 1617.000 ;
    RECT 150.500 1.400 151.340 1617.000 ;
    RECT 151.620 1.400 152.460 1617.000 ;
    RECT 152.740 1.400 153.580 1617.000 ;
    RECT 153.860 1.400 154.700 1617.000 ;
    RECT 154.980 1.400 155.820 1617.000 ;
    RECT 156.100 1.400 156.940 1617.000 ;
    RECT 157.220 1.400 158.060 1617.000 ;
    RECT 158.340 1.400 159.180 1617.000 ;
    RECT 159.460 1.400 160.300 1617.000 ;
    RECT 160.580 1.400 161.420 1617.000 ;
    RECT 161.700 1.400 162.540 1617.000 ;
    RECT 162.820 1.400 163.660 1617.000 ;
    RECT 163.940 1.400 164.780 1617.000 ;
    RECT 165.060 1.400 165.900 1617.000 ;
    RECT 166.180 1.400 167.020 1617.000 ;
    RECT 167.300 1.400 168.140 1617.000 ;
    RECT 168.420 1.400 169.260 1617.000 ;
    RECT 169.540 1.400 170.380 1617.000 ;
    RECT 170.660 1.400 171.500 1617.000 ;
    RECT 171.780 1.400 172.620 1617.000 ;
    RECT 172.900 1.400 173.740 1617.000 ;
    RECT 174.020 1.400 174.860 1617.000 ;
    RECT 175.140 1.400 175.980 1617.000 ;
    RECT 176.260 1.400 177.100 1617.000 ;
    RECT 177.380 1.400 178.220 1617.000 ;
    RECT 178.500 1.400 179.340 1617.000 ;
    RECT 179.620 1.400 180.460 1617.000 ;
    RECT 180.740 1.400 181.580 1617.000 ;
    RECT 181.860 1.400 182.700 1617.000 ;
    RECT 182.980 1.400 183.820 1617.000 ;
    RECT 184.100 1.400 184.940 1617.000 ;
    RECT 185.220 1.400 186.060 1617.000 ;
    RECT 186.340 1.400 187.180 1617.000 ;
    RECT 187.460 1.400 188.300 1617.000 ;
    RECT 188.580 1.400 189.420 1617.000 ;
    RECT 189.700 1.400 190.540 1617.000 ;
    RECT 190.820 1.400 191.660 1617.000 ;
    RECT 191.940 1.400 192.780 1617.000 ;
    RECT 193.060 1.400 193.900 1617.000 ;
    RECT 194.180 1.400 195.020 1617.000 ;
    RECT 195.300 1.400 196.140 1617.000 ;
    RECT 196.420 1.400 197.260 1617.000 ;
    RECT 197.540 1.400 198.380 1617.000 ;
    RECT 198.660 1.400 199.500 1617.000 ;
    RECT 199.780 1.400 200.620 1617.000 ;
    RECT 200.900 1.400 201.740 1617.000 ;
    RECT 202.020 1.400 202.860 1617.000 ;
    RECT 203.140 1.400 203.980 1617.000 ;
    RECT 204.260 1.400 205.100 1617.000 ;
    RECT 205.380 1.400 206.220 1617.000 ;
    RECT 206.500 1.400 207.340 1617.000 ;
    RECT 207.620 1.400 208.460 1617.000 ;
    RECT 208.740 1.400 209.580 1617.000 ;
    RECT 209.860 1.400 210.700 1617.000 ;
    RECT 210.980 1.400 211.820 1617.000 ;
    RECT 212.100 1.400 212.940 1617.000 ;
    RECT 213.220 1.400 214.060 1617.000 ;
    RECT 214.340 1.400 215.180 1617.000 ;
    RECT 215.460 1.400 216.300 1617.000 ;
    RECT 216.580 1.400 217.420 1617.000 ;
    RECT 217.700 1.400 218.540 1617.000 ;
    RECT 218.820 1.400 219.660 1617.000 ;
    RECT 219.940 1.400 220.780 1617.000 ;
    RECT 221.060 1.400 221.900 1617.000 ;
    RECT 222.180 1.400 223.020 1617.000 ;
    RECT 223.300 1.400 224.140 1617.000 ;
    RECT 224.420 1.400 225.260 1617.000 ;
    RECT 225.540 1.400 226.380 1617.000 ;
    RECT 226.660 1.400 227.500 1617.000 ;
    RECT 227.780 1.400 228.620 1617.000 ;
    RECT 228.900 1.400 229.740 1617.000 ;
    RECT 230.020 1.400 230.860 1617.000 ;
    RECT 231.140 1.400 231.980 1617.000 ;
    RECT 232.260 1.400 233.100 1617.000 ;
    RECT 233.380 1.400 234.220 1617.000 ;
    RECT 234.500 1.400 235.340 1617.000 ;
    RECT 235.620 1.400 236.460 1617.000 ;
    RECT 236.740 1.400 237.580 1617.000 ;
    RECT 237.860 1.400 238.700 1617.000 ;
    RECT 238.980 1.400 239.820 1617.000 ;
    RECT 240.100 1.400 240.940 1617.000 ;
    RECT 241.220 1.400 242.060 1617.000 ;
    RECT 242.340 1.400 243.180 1617.000 ;
    RECT 243.460 1.400 244.300 1617.000 ;
    RECT 244.580 1.400 245.420 1617.000 ;
    RECT 245.700 1.400 246.540 1617.000 ;
    RECT 246.820 1.400 247.660 1617.000 ;
    RECT 247.940 1.400 248.780 1617.000 ;
    RECT 249.060 1.400 249.900 1617.000 ;
    RECT 250.180 1.400 251.020 1617.000 ;
    RECT 251.300 1.400 252.140 1617.000 ;
    RECT 252.420 1.400 253.260 1617.000 ;
    RECT 253.540 1.400 254.380 1617.000 ;
    RECT 254.660 1.400 255.500 1617.000 ;
    RECT 255.780 1.400 256.620 1617.000 ;
    RECT 256.900 1.400 257.740 1617.000 ;
    RECT 258.020 1.400 258.860 1617.000 ;
    RECT 259.140 1.400 259.980 1617.000 ;
    RECT 260.260 1.400 261.100 1617.000 ;
    RECT 261.380 1.400 262.220 1617.000 ;
    RECT 262.500 1.400 263.340 1617.000 ;
    RECT 263.620 1.400 264.460 1617.000 ;
    RECT 264.740 1.400 265.580 1617.000 ;
    RECT 265.860 1.400 266.700 1617.000 ;
    RECT 266.980 1.400 267.820 1617.000 ;
    RECT 268.100 1.400 268.940 1617.000 ;
    RECT 269.220 1.400 270.060 1617.000 ;
    RECT 270.340 1.400 271.180 1617.000 ;
    RECT 271.460 1.400 272.300 1617.000 ;
    RECT 272.580 1.400 273.420 1617.000 ;
    RECT 273.700 1.400 274.540 1617.000 ;
    RECT 274.820 1.400 275.660 1617.000 ;
    RECT 275.940 1.400 276.780 1617.000 ;
    RECT 277.060 1.400 277.900 1617.000 ;
    RECT 278.180 1.400 279.020 1617.000 ;
    RECT 279.300 1.400 280.140 1617.000 ;
    RECT 280.420 1.400 281.260 1617.000 ;
    RECT 281.540 1.400 282.380 1617.000 ;
    RECT 282.660 1.400 283.500 1617.000 ;
    RECT 283.780 1.400 284.620 1617.000 ;
    RECT 284.900 1.400 285.740 1617.000 ;
    RECT 286.020 1.400 286.860 1617.000 ;
    RECT 287.140 1.400 287.980 1617.000 ;
    RECT 288.260 1.400 289.100 1617.000 ;
    RECT 289.380 1.400 290.220 1617.000 ;
    RECT 290.500 1.400 291.340 1617.000 ;
    RECT 291.620 1.400 292.460 1617.000 ;
    RECT 292.740 1.400 293.580 1617.000 ;
    RECT 293.860 1.400 294.700 1617.000 ;
    RECT 294.980 1.400 295.820 1617.000 ;
    RECT 296.100 1.400 296.940 1617.000 ;
    RECT 297.220 1.400 298.060 1617.000 ;
    RECT 298.340 1.400 299.180 1617.000 ;
    RECT 299.460 1.400 300.300 1617.000 ;
    RECT 300.580 1.400 301.420 1617.000 ;
    RECT 301.700 1.400 302.540 1617.000 ;
    RECT 302.820 1.400 303.660 1617.000 ;
    RECT 303.940 1.400 304.780 1617.000 ;
    RECT 305.060 1.400 305.900 1617.000 ;
    RECT 306.180 1.400 307.020 1617.000 ;
    RECT 307.300 1.400 308.140 1617.000 ;
    RECT 308.420 1.400 309.260 1617.000 ;
    RECT 309.540 1.400 310.380 1617.000 ;
    RECT 310.660 1.400 311.500 1617.000 ;
    RECT 311.780 1.400 312.620 1617.000 ;
    RECT 312.900 1.400 313.740 1617.000 ;
    RECT 314.020 1.400 314.860 1617.000 ;
    RECT 315.140 1.400 315.980 1617.000 ;
    RECT 316.260 1.400 317.100 1617.000 ;
    RECT 317.380 1.400 318.220 1617.000 ;
    RECT 318.500 1.400 319.340 1617.000 ;
    RECT 319.620 1.400 320.460 1617.000 ;
    RECT 320.740 1.400 321.580 1617.000 ;
    RECT 321.860 1.400 322.700 1617.000 ;
    RECT 322.980 1.400 323.820 1617.000 ;
    RECT 324.100 1.400 324.940 1617.000 ;
    RECT 325.220 1.400 326.060 1617.000 ;
    RECT 326.340 1.400 327.180 1617.000 ;
    RECT 327.460 1.400 328.300 1617.000 ;
    RECT 328.580 1.400 329.420 1617.000 ;
    RECT 329.700 1.400 330.540 1617.000 ;
    RECT 330.820 1.400 331.660 1617.000 ;
    RECT 331.940 1.400 332.780 1617.000 ;
    RECT 333.060 1.400 333.900 1617.000 ;
    RECT 334.180 1.400 335.020 1617.000 ;
    RECT 335.300 1.400 336.140 1617.000 ;
    RECT 336.420 1.400 337.260 1617.000 ;
    RECT 337.540 1.400 338.380 1617.000 ;
    RECT 338.660 1.400 339.500 1617.000 ;
    RECT 339.780 1.400 340.620 1617.000 ;
    RECT 340.900 1.400 341.740 1617.000 ;
    RECT 342.020 1.400 342.860 1617.000 ;
    RECT 343.140 1.400 343.980 1617.000 ;
    RECT 344.260 1.400 345.100 1617.000 ;
    RECT 345.380 1.400 346.220 1617.000 ;
    RECT 346.500 1.400 347.340 1617.000 ;
    RECT 347.620 1.400 348.460 1617.000 ;
    RECT 348.740 1.400 349.580 1617.000 ;
    RECT 349.860 1.400 350.700 1617.000 ;
    RECT 350.980 1.400 351.820 1617.000 ;
    RECT 352.100 1.400 352.940 1617.000 ;
    RECT 353.220 1.400 354.060 1617.000 ;
    RECT 354.340 1.400 355.180 1617.000 ;
    RECT 355.460 1.400 356.300 1617.000 ;
    RECT 356.580 1.400 357.420 1617.000 ;
    RECT 357.700 1.400 358.540 1617.000 ;
    RECT 358.820 1.400 359.660 1617.000 ;
    RECT 359.940 1.400 360.780 1617.000 ;
    RECT 361.060 1.400 361.900 1617.000 ;
    RECT 362.180 1.400 363.020 1617.000 ;
    RECT 363.300 1.400 364.140 1617.000 ;
    RECT 364.420 1.400 365.260 1617.000 ;
    RECT 365.540 1.400 366.380 1617.000 ;
    RECT 366.660 1.400 367.500 1617.000 ;
    RECT 367.780 1.400 368.620 1617.000 ;
    RECT 368.900 1.400 369.740 1617.000 ;
    RECT 370.020 1.400 370.860 1617.000 ;
    RECT 371.140 1.400 371.980 1617.000 ;
    RECT 372.260 1.400 373.100 1617.000 ;
    RECT 373.380 1.400 374.220 1617.000 ;
    RECT 374.500 1.400 375.340 1617.000 ;
    RECT 375.620 1.400 376.460 1617.000 ;
    RECT 376.740 1.400 377.580 1617.000 ;
    RECT 377.860 1.400 378.700 1617.000 ;
    RECT 378.980 1.400 379.820 1617.000 ;
    RECT 380.100 1.400 380.940 1617.000 ;
    RECT 381.220 1.400 382.060 1617.000 ;
    RECT 382.340 1.400 383.180 1617.000 ;
    RECT 383.460 1.400 384.300 1617.000 ;
    RECT 384.580 1.400 385.420 1617.000 ;
    RECT 385.700 1.400 386.540 1617.000 ;
    RECT 386.820 1.400 387.660 1617.000 ;
    RECT 387.940 1.400 388.780 1617.000 ;
    RECT 389.060 1.400 389.900 1617.000 ;
    RECT 390.180 1.400 391.020 1617.000 ;
    RECT 391.300 1.400 392.140 1617.000 ;
    RECT 392.420 1.400 393.260 1617.000 ;
    RECT 393.540 1.400 394.380 1617.000 ;
    RECT 394.660 1.400 395.500 1617.000 ;
    RECT 395.780 1.400 396.620 1617.000 ;
    RECT 396.900 1.400 397.740 1617.000 ;
    RECT 398.020 1.400 398.860 1617.000 ;
    RECT 399.140 1.400 399.980 1617.000 ;
    RECT 400.260 1.400 401.100 1617.000 ;
    RECT 401.380 1.400 402.220 1617.000 ;
    RECT 402.500 1.400 403.340 1617.000 ;
    RECT 403.620 1.400 404.460 1617.000 ;
    RECT 404.740 1.400 405.580 1617.000 ;
    RECT 405.860 1.400 406.700 1617.000 ;
    RECT 406.980 1.400 407.820 1617.000 ;
    RECT 408.100 1.400 408.940 1617.000 ;
    RECT 409.220 1.400 410.060 1617.000 ;
    RECT 410.340 1.400 411.180 1617.000 ;
    RECT 411.460 1.400 412.300 1617.000 ;
    RECT 412.580 1.400 413.420 1617.000 ;
    RECT 413.700 1.400 414.540 1617.000 ;
    RECT 414.820 1.400 415.660 1617.000 ;
    RECT 415.940 1.400 416.780 1617.000 ;
    RECT 417.060 1.400 417.900 1617.000 ;
    RECT 418.180 1.400 419.020 1617.000 ;
    RECT 419.300 1.400 420.140 1617.000 ;
    RECT 420.420 1.400 421.260 1617.000 ;
    RECT 421.540 1.400 422.380 1617.000 ;
    RECT 422.660 1.400 423.500 1617.000 ;
    RECT 423.780 1.400 424.620 1617.000 ;
    RECT 424.900 1.400 425.740 1617.000 ;
    RECT 426.020 1.400 426.860 1617.000 ;
    RECT 427.140 1.400 427.980 1617.000 ;
    RECT 428.260 1.400 429.100 1617.000 ;
    RECT 429.380 1.400 430.220 1617.000 ;
    RECT 430.500 1.400 431.340 1617.000 ;
    RECT 431.620 1.400 432.460 1617.000 ;
    RECT 432.740 1.400 433.580 1617.000 ;
    RECT 433.860 1.400 434.700 1617.000 ;
    RECT 434.980 1.400 435.820 1617.000 ;
    RECT 436.100 1.400 436.940 1617.000 ;
    RECT 437.220 1.400 438.060 1617.000 ;
    RECT 438.340 1.400 439.180 1617.000 ;
    RECT 439.460 1.400 440.300 1617.000 ;
    RECT 440.580 1.400 441.420 1617.000 ;
    RECT 441.700 1.400 442.540 1617.000 ;
    RECT 442.820 1.400 443.660 1617.000 ;
    RECT 443.940 1.400 444.780 1617.000 ;
    RECT 445.060 1.400 445.900 1617.000 ;
    RECT 446.180 1.400 447.020 1617.000 ;
    RECT 447.300 1.400 448.140 1617.000 ;
    RECT 448.420 1.400 449.260 1617.000 ;
    RECT 449.540 1.400 450.380 1617.000 ;
    RECT 450.660 1.400 451.500 1617.000 ;
    RECT 451.780 1.400 452.620 1617.000 ;
    RECT 452.900 1.400 453.740 1617.000 ;
    RECT 454.020 1.400 454.860 1617.000 ;
    RECT 455.140 1.400 455.980 1617.000 ;
    RECT 456.260 1.400 457.100 1617.000 ;
    RECT 457.380 1.400 458.220 1617.000 ;
    RECT 458.500 1.400 459.340 1617.000 ;
    RECT 459.620 1.400 460.460 1617.000 ;
    RECT 460.740 1.400 461.580 1617.000 ;
    RECT 461.860 1.400 462.700 1617.000 ;
    RECT 462.980 1.400 463.820 1617.000 ;
    RECT 464.100 1.400 464.940 1617.000 ;
    RECT 465.220 1.400 466.060 1617.000 ;
    RECT 466.340 1.400 467.180 1617.000 ;
    RECT 467.460 1.400 468.300 1617.000 ;
    RECT 468.580 1.400 469.420 1617.000 ;
    RECT 469.700 1.400 470.540 1617.000 ;
    RECT 470.820 1.400 471.660 1617.000 ;
    RECT 471.940 1.400 472.780 1617.000 ;
    RECT 473.060 1.400 473.900 1617.000 ;
    RECT 474.180 1.400 475.020 1617.000 ;
    RECT 475.300 1.400 476.140 1617.000 ;
    RECT 476.420 1.400 477.260 1617.000 ;
    RECT 477.540 1.400 478.380 1617.000 ;
    RECT 478.660 1.400 479.500 1617.000 ;
    RECT 479.780 1.400 480.620 1617.000 ;
    RECT 480.900 1.400 481.740 1617.000 ;
    RECT 482.020 1.400 482.860 1617.000 ;
    RECT 483.140 1.400 483.980 1617.000 ;
    RECT 484.260 1.400 485.100 1617.000 ;
    RECT 485.380 1.400 486.220 1617.000 ;
    RECT 486.500 1.400 487.340 1617.000 ;
    RECT 487.620 1.400 488.460 1617.000 ;
    RECT 488.740 1.400 489.580 1617.000 ;
    RECT 489.860 1.400 490.700 1617.000 ;
    RECT 490.980 1.400 491.820 1617.000 ;
    RECT 492.100 1.400 492.940 1617.000 ;
    RECT 493.220 1.400 494.060 1617.000 ;
    RECT 494.340 1.400 495.180 1617.000 ;
    RECT 495.460 1.400 496.300 1617.000 ;
    RECT 496.580 1.400 497.420 1617.000 ;
    RECT 497.700 1.400 498.540 1617.000 ;
    RECT 498.820 1.400 499.660 1617.000 ;
    RECT 499.940 1.400 500.780 1617.000 ;
    RECT 501.060 1.400 501.900 1617.000 ;
    RECT 502.180 1.400 503.020 1617.000 ;
    RECT 503.300 1.400 504.140 1617.000 ;
    RECT 504.420 1.400 505.260 1617.000 ;
    RECT 505.540 1.400 506.380 1617.000 ;
    RECT 506.660 1.400 507.500 1617.000 ;
    RECT 507.780 1.400 508.620 1617.000 ;
    RECT 508.900 1.400 509.740 1617.000 ;
    RECT 510.020 1.400 510.860 1617.000 ;
    RECT 511.140 1.400 511.980 1617.000 ;
    RECT 512.260 1.400 513.100 1617.000 ;
    RECT 513.380 1.400 514.220 1617.000 ;
    RECT 514.500 1.400 515.340 1617.000 ;
    RECT 515.620 1.400 516.460 1617.000 ;
    RECT 516.740 1.400 517.580 1617.000 ;
    RECT 517.860 1.400 518.700 1617.000 ;
    RECT 518.980 1.400 519.820 1617.000 ;
    RECT 520.100 1.400 520.940 1617.000 ;
    RECT 521.220 1.400 522.060 1617.000 ;
    RECT 522.340 1.400 523.180 1617.000 ;
    RECT 523.460 1.400 524.300 1617.000 ;
    RECT 524.580 1.400 525.420 1617.000 ;
    RECT 525.700 1.400 526.540 1617.000 ;
    RECT 526.820 1.400 527.660 1617.000 ;
    RECT 527.940 1.400 528.780 1617.000 ;
    RECT 529.060 1.400 529.900 1617.000 ;
    RECT 530.180 1.400 531.020 1617.000 ;
    RECT 531.300 1.400 532.140 1617.000 ;
    RECT 532.420 1.400 533.260 1617.000 ;
    RECT 533.540 1.400 534.380 1617.000 ;
    RECT 534.660 1.400 535.500 1617.000 ;
    RECT 535.780 1.400 536.620 1617.000 ;
    RECT 536.900 1.400 537.740 1617.000 ;
    RECT 538.020 1.400 538.860 1617.000 ;
    RECT 539.140 1.400 539.980 1617.000 ;
    RECT 540.260 1.400 541.100 1617.000 ;
    RECT 541.380 1.400 542.220 1617.000 ;
    RECT 542.500 1.400 543.340 1617.000 ;
    RECT 543.620 1.400 544.460 1617.000 ;
    RECT 544.740 1.400 545.580 1617.000 ;
    RECT 545.860 1.400 546.700 1617.000 ;
    RECT 546.980 1.400 547.820 1617.000 ;
    RECT 548.100 1.400 548.940 1617.000 ;
    RECT 549.220 1.400 550.060 1617.000 ;
    RECT 550.340 1.400 551.180 1617.000 ;
    RECT 551.460 1.400 552.300 1617.000 ;
    RECT 552.580 1.400 553.420 1617.000 ;
    RECT 553.700 1.400 554.540 1617.000 ;
    RECT 554.820 1.400 555.660 1617.000 ;
    RECT 555.940 1.400 556.780 1617.000 ;
    RECT 557.060 1.400 557.900 1617.000 ;
    RECT 558.180 1.400 559.020 1617.000 ;
    RECT 559.300 1.400 560.140 1617.000 ;
    RECT 560.420 1.400 561.260 1617.000 ;
    RECT 561.540 1.400 562.380 1617.000 ;
    RECT 562.660 1.400 563.500 1617.000 ;
    RECT 563.780 1.400 564.620 1617.000 ;
    RECT 564.900 1.400 565.740 1617.000 ;
    RECT 566.020 1.400 566.860 1617.000 ;
    RECT 567.140 1.400 567.980 1617.000 ;
    RECT 568.260 1.400 569.100 1617.000 ;
    RECT 569.380 1.400 570.220 1617.000 ;
    RECT 570.500 1.400 571.340 1617.000 ;
    RECT 571.620 1.400 572.460 1617.000 ;
    RECT 572.740 1.400 573.580 1617.000 ;
    RECT 573.860 1.400 574.700 1617.000 ;
    RECT 574.980 1.400 575.820 1617.000 ;
    RECT 576.100 1.400 576.940 1617.000 ;
    RECT 577.220 1.400 578.060 1617.000 ;
    RECT 578.340 1.400 579.180 1617.000 ;
    RECT 579.460 1.400 580.300 1617.000 ;
    RECT 580.580 1.400 581.420 1617.000 ;
    RECT 581.700 1.400 582.540 1617.000 ;
    RECT 582.820 1.400 583.660 1617.000 ;
    RECT 583.940 1.400 584.780 1617.000 ;
    RECT 585.060 1.400 585.900 1617.000 ;
    RECT 586.180 1.400 587.020 1617.000 ;
    RECT 587.300 1.400 588.140 1617.000 ;
    RECT 588.420 1.400 589.260 1617.000 ;
    RECT 589.540 1.400 590.380 1617.000 ;
    RECT 590.660 1.400 591.500 1617.000 ;
    RECT 591.780 1.400 592.620 1617.000 ;
    RECT 592.900 1.400 593.740 1617.000 ;
    RECT 594.020 1.400 594.860 1617.000 ;
    RECT 595.140 1.400 595.980 1617.000 ;
    RECT 596.260 1.400 597.100 1617.000 ;
    RECT 597.380 1.400 598.220 1617.000 ;
    RECT 598.500 1.400 599.340 1617.000 ;
    RECT 599.620 1.400 600.460 1617.000 ;
    RECT 600.740 1.400 601.580 1617.000 ;
    RECT 601.860 1.400 602.700 1617.000 ;
    RECT 602.980 1.400 603.820 1617.000 ;
    RECT 604.100 1.400 604.940 1617.000 ;
    RECT 605.220 1.400 606.060 1617.000 ;
    RECT 606.340 1.400 607.180 1617.000 ;
    RECT 607.460 1.400 608.300 1617.000 ;
    RECT 608.580 1.400 609.420 1617.000 ;
    RECT 609.700 1.400 610.540 1617.000 ;
    RECT 610.820 1.400 611.660 1617.000 ;
    RECT 611.940 1.400 612.780 1617.000 ;
    RECT 613.060 1.400 613.900 1617.000 ;
    RECT 614.180 1.400 615.020 1617.000 ;
    RECT 615.300 1.400 616.140 1617.000 ;
    RECT 616.420 1.400 617.260 1617.000 ;
    RECT 617.540 1.400 618.380 1617.000 ;
    RECT 618.660 1.400 619.500 1617.000 ;
    RECT 619.780 1.400 620.620 1617.000 ;
    RECT 620.900 1.400 621.740 1617.000 ;
    RECT 622.020 1.400 622.860 1617.000 ;
    RECT 623.140 1.400 623.980 1617.000 ;
    RECT 624.260 1.400 625.100 1617.000 ;
    RECT 625.380 1.400 626.220 1617.000 ;
    RECT 626.500 1.400 627.340 1617.000 ;
    RECT 627.620 1.400 628.460 1617.000 ;
    RECT 628.740 1.400 629.580 1617.000 ;
    RECT 629.860 1.400 630.700 1617.000 ;
    RECT 630.980 1.400 631.820 1617.000 ;
    RECT 632.100 1.400 632.940 1617.000 ;
    RECT 633.220 1.400 634.060 1617.000 ;
    RECT 634.340 1.400 635.180 1617.000 ;
    RECT 635.460 1.400 636.300 1617.000 ;
    RECT 636.580 1.400 637.420 1617.000 ;
    RECT 637.700 1.400 638.540 1617.000 ;
    RECT 638.820 1.400 639.660 1617.000 ;
    RECT 639.940 1.400 640.780 1617.000 ;
    RECT 641.060 1.400 641.900 1617.000 ;
    RECT 642.180 1.400 643.020 1617.000 ;
    RECT 643.300 1.400 644.140 1617.000 ;
    RECT 644.420 1.400 645.260 1617.000 ;
    RECT 645.540 1.400 646.380 1617.000 ;
    RECT 646.660 1.400 647.500 1617.000 ;
    RECT 647.780 1.400 648.620 1617.000 ;
    RECT 648.900 1.400 649.740 1617.000 ;
    RECT 650.020 1.400 650.860 1617.000 ;
    RECT 651.140 1.400 651.980 1617.000 ;
    RECT 652.260 1.400 653.100 1617.000 ;
    RECT 653.380 1.400 654.220 1617.000 ;
    RECT 654.500 1.400 655.340 1617.000 ;
    RECT 655.620 1.400 656.460 1617.000 ;
    RECT 656.740 1.400 657.580 1617.000 ;
    RECT 657.860 1.400 658.700 1617.000 ;
    RECT 658.980 1.400 659.820 1617.000 ;
    RECT 660.100 1.400 660.940 1617.000 ;
    RECT 661.220 1.400 662.060 1617.000 ;
    RECT 662.340 1.400 663.180 1617.000 ;
    RECT 663.460 1.400 664.300 1617.000 ;
    RECT 664.580 1.400 665.420 1617.000 ;
    RECT 665.700 1.400 666.540 1617.000 ;
    RECT 666.820 1.400 667.660 1617.000 ;
    RECT 667.940 1.400 668.780 1617.000 ;
    RECT 669.060 1.400 669.900 1617.000 ;
    RECT 670.180 1.400 671.020 1617.000 ;
    RECT 671.300 1.400 672.140 1617.000 ;
    RECT 672.420 1.400 673.260 1617.000 ;
    RECT 673.540 1.400 674.380 1617.000 ;
    RECT 674.660 1.400 675.500 1617.000 ;
    RECT 675.780 1.400 676.620 1617.000 ;
    RECT 676.900 1.400 677.740 1617.000 ;
    RECT 678.020 1.400 678.860 1617.000 ;
    RECT 679.140 1.400 679.980 1617.000 ;
    RECT 680.260 1.400 681.100 1617.000 ;
    RECT 681.380 1.400 682.220 1617.000 ;
    RECT 682.500 1.400 683.340 1617.000 ;
    RECT 683.620 1.400 684.460 1617.000 ;
    RECT 684.740 1.400 685.580 1617.000 ;
    RECT 685.860 1.400 686.700 1617.000 ;
    RECT 686.980 1.400 687.820 1617.000 ;
    RECT 688.100 1.400 688.940 1617.000 ;
    RECT 689.220 1.400 690.060 1617.000 ;
    RECT 690.340 1.400 691.180 1617.000 ;
    RECT 691.460 1.400 692.300 1617.000 ;
    RECT 692.580 1.400 693.420 1617.000 ;
    RECT 693.700 1.400 694.540 1617.000 ;
    RECT 694.820 1.400 695.660 1617.000 ;
    RECT 695.940 1.400 696.780 1617.000 ;
    RECT 697.060 1.400 697.900 1617.000 ;
    RECT 698.180 1.400 699.020 1617.000 ;
    RECT 699.300 1.400 700.140 1617.000 ;
    RECT 700.420 1.400 701.260 1617.000 ;
    RECT 701.540 1.400 702.380 1617.000 ;
    RECT 702.660 1.400 703.500 1617.000 ;
    RECT 703.780 1.400 704.620 1617.000 ;
    RECT 704.900 1.400 705.740 1617.000 ;
    RECT 706.020 1.400 706.860 1617.000 ;
    RECT 707.140 1.400 707.980 1617.000 ;
    RECT 708.260 1.400 709.100 1617.000 ;
    RECT 709.380 1.400 710.220 1617.000 ;
    RECT 710.500 1.400 711.340 1617.000 ;
    RECT 711.620 1.400 712.460 1617.000 ;
    RECT 712.740 1.400 713.580 1617.000 ;
    RECT 713.860 1.400 714.700 1617.000 ;
    RECT 714.980 1.400 715.820 1617.000 ;
    RECT 716.100 1.400 716.940 1617.000 ;
    RECT 717.220 1.400 718.060 1617.000 ;
    RECT 718.340 1.400 719.180 1617.000 ;
    RECT 719.460 1.400 720.300 1617.000 ;
    RECT 720.580 1.400 721.420 1617.000 ;
    RECT 721.700 1.400 722.540 1617.000 ;
    RECT 722.820 1.400 723.660 1617.000 ;
    RECT 723.940 1.400 724.780 1617.000 ;
    RECT 725.060 1.400 725.900 1617.000 ;
    RECT 726.180 1.400 727.020 1617.000 ;
    RECT 727.300 1.400 728.140 1617.000 ;
    RECT 728.420 1.400 729.260 1617.000 ;
    RECT 729.540 1.400 730.380 1617.000 ;
    RECT 730.660 1.400 731.500 1617.000 ;
    RECT 731.780 1.400 732.620 1617.000 ;
    RECT 732.900 1.400 733.740 1617.000 ;
    RECT 734.020 1.400 734.860 1617.000 ;
    RECT 735.140 1.400 735.980 1617.000 ;
    RECT 736.260 1.400 737.100 1617.000 ;
    RECT 737.380 1.400 738.220 1617.000 ;
    RECT 738.500 1.400 739.340 1617.000 ;
    RECT 739.620 1.400 740.460 1617.000 ;
    RECT 740.740 1.400 741.580 1617.000 ;
    RECT 741.860 1.400 742.700 1617.000 ;
    RECT 742.980 1.400 743.820 1617.000 ;
    RECT 744.100 1.400 744.940 1617.000 ;
    RECT 745.220 1.400 746.060 1617.000 ;
    RECT 746.340 1.400 747.180 1617.000 ;
    RECT 747.460 1.400 748.300 1617.000 ;
    RECT 748.580 1.400 749.420 1617.000 ;
    RECT 749.700 1.400 750.540 1617.000 ;
    RECT 750.820 1.400 751.660 1617.000 ;
    RECT 751.940 1.400 752.780 1617.000 ;
    RECT 753.060 1.400 753.900 1617.000 ;
    RECT 754.180 1.400 755.020 1617.000 ;
    RECT 755.300 1.400 756.140 1617.000 ;
    RECT 756.420 1.400 757.260 1617.000 ;
    RECT 757.540 1.400 758.380 1617.000 ;
    RECT 758.660 1.400 759.500 1617.000 ;
    RECT 759.780 1.400 760.620 1617.000 ;
    RECT 760.900 1.400 761.740 1617.000 ;
    RECT 762.020 1.400 762.860 1617.000 ;
    RECT 763.140 1.400 763.980 1617.000 ;
    RECT 764.260 1.400 765.100 1617.000 ;
    RECT 765.380 1.400 766.220 1617.000 ;
    RECT 766.500 1.400 767.340 1617.000 ;
    RECT 767.620 1.400 768.460 1617.000 ;
    RECT 768.740 1.400 769.580 1617.000 ;
    RECT 769.860 1.400 770.700 1617.000 ;
    RECT 770.980 1.400 771.820 1617.000 ;
    RECT 772.100 1.400 772.940 1617.000 ;
    RECT 773.220 1.400 774.060 1617.000 ;
    RECT 774.340 1.400 775.180 1617.000 ;
    RECT 775.460 1.400 776.300 1617.000 ;
    RECT 776.580 1.400 777.420 1617.000 ;
    RECT 777.700 1.400 778.540 1617.000 ;
    RECT 778.820 1.400 779.660 1617.000 ;
    RECT 779.940 1.400 780.780 1617.000 ;
    RECT 781.060 1.400 781.900 1617.000 ;
    RECT 782.180 1.400 783.020 1617.000 ;
    RECT 783.300 1.400 784.140 1617.000 ;
    RECT 784.420 1.400 785.260 1617.000 ;
    RECT 785.540 1.400 786.380 1617.000 ;
    RECT 786.660 1.400 787.500 1617.000 ;
    RECT 787.780 1.400 788.620 1617.000 ;
    RECT 788.900 1.400 789.740 1617.000 ;
    RECT 790.020 1.400 790.860 1617.000 ;
    RECT 791.140 1.400 791.980 1617.000 ;
    RECT 792.260 1.400 793.100 1617.000 ;
    RECT 793.380 1.400 794.220 1617.000 ;
    RECT 794.500 1.400 795.340 1617.000 ;
    RECT 795.620 1.400 796.460 1617.000 ;
    RECT 796.740 1.400 797.580 1617.000 ;
    RECT 797.860 1.400 798.700 1617.000 ;
    RECT 798.980 1.400 799.820 1617.000 ;
    RECT 800.100 1.400 800.940 1617.000 ;
    RECT 801.220 1.400 802.060 1617.000 ;
    RECT 802.340 1.400 803.180 1617.000 ;
    RECT 803.460 1.400 804.300 1617.000 ;
    RECT 804.580 1.400 805.420 1617.000 ;
    RECT 805.700 1.400 806.540 1617.000 ;
    RECT 806.820 1.400 807.660 1617.000 ;
    RECT 807.940 1.400 808.780 1617.000 ;
    RECT 809.060 1.400 809.900 1617.000 ;
    RECT 810.180 1.400 811.020 1617.000 ;
    RECT 811.300 1.400 812.140 1617.000 ;
    RECT 812.420 1.400 813.260 1617.000 ;
    RECT 813.540 1.400 814.380 1617.000 ;
    RECT 814.660 1.400 815.500 1617.000 ;
    RECT 815.780 1.400 816.620 1617.000 ;
    RECT 816.900 1.400 817.740 1617.000 ;
    RECT 818.020 1.400 818.860 1617.000 ;
    RECT 819.140 1.400 819.980 1617.000 ;
    RECT 820.260 1.400 821.100 1617.000 ;
    RECT 821.380 1.400 822.220 1617.000 ;
    RECT 822.500 1.400 823.340 1617.000 ;
    RECT 823.620 1.400 824.460 1617.000 ;
    RECT 824.740 1.400 825.580 1617.000 ;
    RECT 825.860 1.400 826.700 1617.000 ;
    RECT 826.980 1.400 827.820 1617.000 ;
    RECT 828.100 1.400 828.940 1617.000 ;
    RECT 829.220 1.400 830.060 1617.000 ;
    RECT 830.340 1.400 831.180 1617.000 ;
    RECT 831.460 1.400 832.300 1617.000 ;
    RECT 832.580 1.400 833.420 1617.000 ;
    RECT 833.700 1.400 834.540 1617.000 ;
    RECT 834.820 1.400 835.660 1617.000 ;
    RECT 835.940 1.400 836.780 1617.000 ;
    RECT 837.060 1.400 837.900 1617.000 ;
    RECT 838.180 1.400 839.020 1617.000 ;
    RECT 839.300 1.400 840.140 1617.000 ;
    RECT 840.420 1.400 841.260 1617.000 ;
    RECT 841.540 1.400 842.380 1617.000 ;
    RECT 842.660 1.400 843.500 1617.000 ;
    RECT 843.780 1.400 844.620 1617.000 ;
    RECT 844.900 1.400 845.740 1617.000 ;
    RECT 846.020 1.400 846.860 1617.000 ;
    RECT 847.140 1.400 847.980 1617.000 ;
    RECT 848.260 1.400 849.100 1617.000 ;
    RECT 849.380 1.400 850.220 1617.000 ;
    RECT 850.500 1.400 851.340 1617.000 ;
    RECT 851.620 1.400 852.460 1617.000 ;
    RECT 852.740 1.400 853.580 1617.000 ;
    RECT 853.860 1.400 854.700 1617.000 ;
    RECT 854.980 1.400 855.820 1617.000 ;
    RECT 856.100 1.400 856.940 1617.000 ;
    RECT 857.220 1.400 858.060 1617.000 ;
    RECT 858.340 1.400 859.180 1617.000 ;
    RECT 859.460 1.400 860.300 1617.000 ;
    RECT 860.580 1.400 861.420 1617.000 ;
    RECT 861.700 1.400 862.540 1617.000 ;
    RECT 862.820 1.400 863.660 1617.000 ;
    RECT 863.940 1.400 864.780 1617.000 ;
    RECT 865.060 1.400 865.900 1617.000 ;
    RECT 866.180 1.400 867.020 1617.000 ;
    RECT 867.300 1.400 868.140 1617.000 ;
    RECT 868.420 1.400 869.260 1617.000 ;
    RECT 869.540 1.400 870.380 1617.000 ;
    RECT 870.660 1.400 871.500 1617.000 ;
    RECT 871.780 1.400 872.620 1617.000 ;
    RECT 872.900 1.400 873.740 1617.000 ;
    RECT 874.020 1.400 874.860 1617.000 ;
    RECT 875.140 1.400 875.980 1617.000 ;
    RECT 876.260 1.400 877.100 1617.000 ;
    RECT 877.380 1.400 878.220 1617.000 ;
    RECT 878.500 1.400 879.340 1617.000 ;
    RECT 879.620 1.400 880.460 1617.000 ;
    RECT 880.740 1.400 881.580 1617.000 ;
    RECT 881.860 1.400 882.700 1617.000 ;
    RECT 882.980 1.400 883.820 1617.000 ;
    RECT 884.100 1.400 884.940 1617.000 ;
    RECT 885.220 1.400 886.060 1617.000 ;
    RECT 886.340 1.400 887.180 1617.000 ;
    RECT 887.460 1.400 888.300 1617.000 ;
    RECT 888.580 1.400 889.420 1617.000 ;
    RECT 889.700 1.400 890.540 1617.000 ;
    RECT 890.820 1.400 891.660 1617.000 ;
    RECT 891.940 1.400 892.780 1617.000 ;
    RECT 893.060 1.400 893.900 1617.000 ;
    RECT 894.180 1.400 895.020 1617.000 ;
    RECT 895.300 1.400 896.140 1617.000 ;
    RECT 896.420 1.400 897.260 1617.000 ;
    RECT 897.540 1.400 898.380 1617.000 ;
    RECT 898.660 1.400 899.500 1617.000 ;
    RECT 899.780 1.400 900.620 1617.000 ;
    RECT 900.900 1.400 901.740 1617.000 ;
    RECT 902.020 1.400 902.860 1617.000 ;
    RECT 903.140 1.400 903.980 1617.000 ;
    RECT 904.260 1.400 905.100 1617.000 ;
    RECT 905.380 1.400 906.220 1617.000 ;
    RECT 906.500 1.400 907.340 1617.000 ;
    RECT 907.620 1.400 908.460 1617.000 ;
    RECT 908.740 1.400 909.580 1617.000 ;
    RECT 909.860 1.400 910.700 1617.000 ;
    RECT 910.980 1.400 911.820 1617.000 ;
    RECT 912.100 1.400 912.940 1617.000 ;
    RECT 913.220 1.400 914.060 1617.000 ;
    RECT 914.340 1.400 915.180 1617.000 ;
    RECT 915.460 1.400 916.300 1617.000 ;
    RECT 916.580 1.400 917.420 1617.000 ;
    RECT 917.700 1.400 918.540 1617.000 ;
    RECT 918.820 1.400 919.660 1617.000 ;
    RECT 919.940 1.400 920.780 1617.000 ;
    RECT 921.060 1.400 921.900 1617.000 ;
    RECT 922.180 1.400 923.020 1617.000 ;
    RECT 923.300 1.400 924.140 1617.000 ;
    RECT 924.420 1.400 925.260 1617.000 ;
    RECT 925.540 1.400 926.380 1617.000 ;
    RECT 926.660 1.400 927.500 1617.000 ;
    RECT 927.780 1.400 928.620 1617.000 ;
    RECT 928.900 1.400 929.740 1617.000 ;
    RECT 930.020 1.400 930.860 1617.000 ;
    RECT 931.140 1.400 931.980 1617.000 ;
    RECT 932.260 1.400 933.100 1617.000 ;
    RECT 933.380 1.400 934.220 1617.000 ;
    RECT 934.500 1.400 935.340 1617.000 ;
    RECT 935.620 1.400 936.460 1617.000 ;
    RECT 936.740 1.400 937.580 1617.000 ;
    RECT 937.860 1.400 938.700 1617.000 ;
    RECT 938.980 1.400 939.820 1617.000 ;
    RECT 940.100 1.400 940.940 1617.000 ;
    RECT 941.220 1.400 942.060 1617.000 ;
    RECT 942.340 1.400 943.180 1617.000 ;
    RECT 943.460 1.400 944.300 1617.000 ;
    RECT 944.580 1.400 945.420 1617.000 ;
    RECT 945.700 1.400 946.540 1617.000 ;
    RECT 946.820 1.400 947.660 1617.000 ;
    RECT 947.940 1.400 948.780 1617.000 ;
    RECT 949.060 1.400 949.900 1617.000 ;
    RECT 950.180 1.400 951.020 1617.000 ;
    RECT 951.300 1.400 952.140 1617.000 ;
    RECT 952.420 1.400 953.260 1617.000 ;
    RECT 953.540 1.400 954.380 1617.000 ;
    RECT 954.660 1.400 955.500 1617.000 ;
    RECT 955.780 1.400 956.620 1617.000 ;
    RECT 956.900 1.400 957.740 1617.000 ;
    RECT 958.020 1.400 958.860 1617.000 ;
    RECT 959.140 1.400 959.980 1617.000 ;
    RECT 960.260 1.400 961.100 1617.000 ;
    RECT 961.380 1.400 962.220 1617.000 ;
    RECT 962.500 1.400 963.340 1617.000 ;
    RECT 963.620 1.400 964.460 1617.000 ;
    RECT 964.740 1.400 965.580 1617.000 ;
    RECT 965.860 1.400 966.700 1617.000 ;
    RECT 966.980 1.400 967.820 1617.000 ;
    RECT 968.100 1.400 968.940 1617.000 ;
    RECT 969.220 1.400 970.060 1617.000 ;
    RECT 970.340 1.400 971.180 1617.000 ;
    RECT 971.460 1.400 972.300 1617.000 ;
    RECT 972.580 1.400 973.420 1617.000 ;
    RECT 973.700 1.400 974.540 1617.000 ;
    RECT 974.820 1.400 975.660 1617.000 ;
    RECT 975.940 1.400 976.780 1617.000 ;
    RECT 977.060 1.400 977.900 1617.000 ;
    RECT 978.180 1.400 979.020 1617.000 ;
    RECT 979.300 1.400 980.140 1617.000 ;
    RECT 980.420 1.400 981.260 1617.000 ;
    RECT 981.540 1.400 982.380 1617.000 ;
    RECT 982.660 1.400 983.500 1617.000 ;
    RECT 983.780 1.400 984.620 1617.000 ;
    RECT 984.900 1.400 985.740 1617.000 ;
    RECT 986.020 1.400 986.860 1617.000 ;
    RECT 987.140 1.400 987.980 1617.000 ;
    RECT 988.260 1.400 989.100 1617.000 ;
    RECT 989.380 1.400 990.220 1617.000 ;
    RECT 990.500 1.400 991.340 1617.000 ;
    RECT 991.620 1.400 992.460 1617.000 ;
    RECT 992.740 1.400 993.580 1617.000 ;
    RECT 993.860 1.400 994.700 1617.000 ;
    RECT 994.980 1.400 995.820 1617.000 ;
    RECT 996.100 1.400 996.940 1617.000 ;
    RECT 997.220 1.400 998.060 1617.000 ;
    RECT 998.340 1.400 999.180 1617.000 ;
    RECT 999.460 1.400 1000.300 1617.000 ;
    RECT 1000.580 1.400 1001.420 1617.000 ;
    RECT 1001.700 1.400 1002.540 1617.000 ;
    RECT 1002.820 1.400 1003.660 1617.000 ;
    RECT 1003.940 1.400 1004.780 1617.000 ;
    RECT 1005.060 1.400 1005.900 1617.000 ;
    RECT 1006.180 1.400 1007.020 1617.000 ;
    RECT 1007.300 1.400 1008.140 1617.000 ;
    RECT 1008.420 1.400 1009.260 1617.000 ;
    RECT 1009.540 1.400 1010.380 1617.000 ;
    RECT 1010.660 1.400 1011.500 1617.000 ;
    RECT 1011.780 1.400 1012.620 1617.000 ;
    RECT 1012.900 1.400 1013.740 1617.000 ;
    RECT 1014.020 1.400 1014.860 1617.000 ;
    RECT 1015.140 1.400 1015.980 1617.000 ;
    RECT 1016.260 1.400 1017.100 1617.000 ;
    RECT 1017.380 1.400 1018.220 1617.000 ;
    RECT 1018.500 1.400 1019.340 1617.000 ;
    RECT 1019.620 1.400 1020.460 1617.000 ;
    RECT 1020.740 1.400 1021.580 1617.000 ;
    RECT 1021.860 1.400 1022.700 1617.000 ;
    RECT 1022.980 1.400 1023.820 1617.000 ;
    RECT 1024.100 1.400 1024.940 1617.000 ;
    RECT 1025.220 1.400 1026.060 1617.000 ;
    RECT 1026.340 1.400 1027.180 1617.000 ;
    RECT 1027.460 1.400 1028.300 1617.000 ;
    RECT 1028.580 1.400 1029.420 1617.000 ;
    RECT 1029.700 1.400 1030.540 1617.000 ;
    RECT 1030.820 1.400 1031.660 1617.000 ;
    RECT 1031.940 1.400 1032.780 1617.000 ;
    RECT 1033.060 1.400 1033.900 1617.000 ;
    RECT 1034.180 1.400 1035.020 1617.000 ;
    RECT 1035.300 1.400 1036.140 1617.000 ;
    RECT 1036.420 1.400 1037.260 1617.000 ;
    RECT 1037.540 1.400 1038.380 1617.000 ;
    RECT 1038.660 1.400 1039.500 1617.000 ;
    RECT 1039.780 1.400 1040.620 1617.000 ;
    RECT 1040.900 1.400 1041.740 1617.000 ;
    RECT 1042.020 1.400 1042.860 1617.000 ;
    RECT 1043.140 1.400 1043.980 1617.000 ;
    RECT 1044.260 1.400 1045.100 1617.000 ;
    RECT 1045.380 1.400 1046.220 1617.000 ;
    RECT 1046.500 1.400 1047.340 1617.000 ;
    RECT 1047.620 1.400 1048.460 1617.000 ;
    RECT 1048.740 1.400 1049.580 1617.000 ;
    RECT 1049.860 1.400 1050.700 1617.000 ;
    RECT 1050.980 1.400 1051.820 1617.000 ;
    RECT 1052.100 1.400 1052.940 1617.000 ;
    RECT 1053.220 1.400 1054.060 1617.000 ;
    RECT 1054.340 1.400 1055.180 1617.000 ;
    RECT 1055.460 1.400 1056.300 1617.000 ;
    RECT 1056.580 1.400 1057.420 1617.000 ;
    RECT 1057.700 1.400 1058.540 1617.000 ;
    RECT 1058.820 1.400 1059.660 1617.000 ;
    RECT 1059.940 1.400 1060.780 1617.000 ;
    RECT 1061.060 1.400 1061.900 1617.000 ;
    RECT 1062.180 1.400 1063.020 1617.000 ;
    RECT 1063.300 1.400 1064.140 1617.000 ;
    RECT 1064.420 1.400 1065.260 1617.000 ;
    RECT 1065.540 1.400 1066.380 1617.000 ;
    RECT 1066.660 1.400 1067.500 1617.000 ;
    RECT 1067.780 1.400 1068.620 1617.000 ;
    RECT 1068.900 1.400 1069.740 1617.000 ;
    RECT 1070.020 1.400 1070.860 1617.000 ;
    RECT 1071.140 1.400 1071.980 1617.000 ;
    RECT 1072.260 1.400 1073.100 1617.000 ;
    RECT 1073.380 1.400 1074.220 1617.000 ;
    RECT 1074.500 1.400 1075.340 1617.000 ;
    RECT 1075.620 1.400 1076.460 1617.000 ;
    RECT 1076.740 1.400 1077.580 1617.000 ;
    RECT 1077.860 1.400 1078.700 1617.000 ;
    RECT 1078.980 1.400 1079.820 1617.000 ;
    RECT 1080.100 1.400 1080.940 1617.000 ;
    RECT 1081.220 1.400 1082.060 1617.000 ;
    RECT 1082.340 1.400 1083.180 1617.000 ;
    RECT 1083.460 1.400 1084.300 1617.000 ;
    RECT 1084.580 1.400 1085.420 1617.000 ;
    RECT 1085.700 1.400 1086.540 1617.000 ;
    RECT 1086.820 1.400 1087.660 1617.000 ;
    RECT 1087.940 1.400 1088.780 1617.000 ;
    RECT 1089.060 1.400 1089.900 1617.000 ;
    RECT 1090.180 1.400 1091.020 1617.000 ;
    RECT 1091.300 1.400 1092.140 1617.000 ;
    RECT 1092.420 1.400 1093.260 1617.000 ;
    RECT 1093.540 1.400 1094.380 1617.000 ;
    RECT 1094.660 1.400 1095.500 1617.000 ;
    RECT 1095.780 1.400 1096.620 1617.000 ;
    RECT 1096.900 1.400 1097.740 1617.000 ;
    RECT 1098.020 1.400 1098.860 1617.000 ;
    RECT 1099.140 1.400 1099.980 1617.000 ;
    RECT 1100.260 1.400 1101.100 1617.000 ;
    RECT 1101.380 1.400 1102.220 1617.000 ;
    RECT 1102.500 1.400 1103.340 1617.000 ;
    RECT 1103.620 1.400 1104.460 1617.000 ;
    RECT 1104.740 1.400 1105.580 1617.000 ;
    RECT 1105.860 1.400 1106.700 1617.000 ;
    RECT 1106.980 1.400 1107.820 1617.000 ;
    RECT 1108.100 1.400 1108.940 1617.000 ;
    RECT 1109.220 1.400 1110.060 1617.000 ;
    RECT 1110.340 1.400 1111.180 1617.000 ;
    RECT 1111.460 1.400 1112.300 1617.000 ;
    RECT 1112.580 1.400 1113.420 1617.000 ;
    RECT 1113.700 1.400 1114.540 1617.000 ;
    RECT 1114.820 1.400 1115.660 1617.000 ;
    RECT 1115.940 1.400 1116.780 1617.000 ;
    RECT 1117.060 1.400 1117.900 1617.000 ;
    RECT 1118.180 1.400 1119.020 1617.000 ;
    RECT 1119.300 1.400 1120.140 1617.000 ;
    RECT 1120.420 1.400 1121.260 1617.000 ;
    RECT 1121.540 1.400 1122.380 1617.000 ;
    RECT 1122.660 1.400 1123.500 1617.000 ;
    RECT 1123.780 1.400 1124.620 1617.000 ;
    RECT 1124.900 1.400 1125.740 1617.000 ;
    RECT 1126.020 1.400 1126.860 1617.000 ;
    RECT 1127.140 1.400 1127.980 1617.000 ;
    RECT 1128.260 1.400 1129.100 1617.000 ;
    RECT 1129.380 1.400 1130.220 1617.000 ;
    RECT 1130.500 1.400 1131.340 1617.000 ;
    RECT 1131.620 1.400 1132.460 1617.000 ;
    RECT 1132.740 1.400 1133.580 1617.000 ;
    RECT 1133.860 1.400 1134.700 1617.000 ;
    RECT 1134.980 1.400 1135.820 1617.000 ;
    RECT 1136.100 1.400 1136.940 1617.000 ;
    RECT 1137.220 1.400 1138.060 1617.000 ;
    RECT 1138.340 1.400 1139.180 1617.000 ;
    RECT 1139.460 1.400 1140.300 1617.000 ;
    RECT 1140.580 1.400 1141.420 1617.000 ;
    RECT 1141.700 1.400 1142.540 1617.000 ;
    RECT 1142.820 1.400 1143.660 1617.000 ;
    RECT 1143.940 1.400 1144.780 1617.000 ;
    RECT 1145.060 1.400 1145.900 1617.000 ;
    RECT 1146.180 1.400 1147.020 1617.000 ;
    RECT 1147.300 1.400 1148.140 1617.000 ;
    RECT 1148.420 1.400 1149.260 1617.000 ;
    RECT 1149.540 1.400 1150.380 1617.000 ;
    RECT 1150.660 1.400 1151.500 1617.000 ;
    RECT 1151.780 1.400 1152.620 1617.000 ;
    RECT 1152.900 1.400 1153.740 1617.000 ;
    RECT 1154.020 1.400 1154.860 1617.000 ;
    RECT 1155.140 1.400 1155.980 1617.000 ;
    RECT 1156.260 1.400 1157.100 1617.000 ;
    RECT 1157.380 1.400 1158.220 1617.000 ;
    RECT 1158.500 1.400 1159.340 1617.000 ;
    RECT 1159.620 1.400 1160.460 1617.000 ;
    RECT 1160.740 1.400 1161.580 1617.000 ;
    RECT 1161.860 1.400 1162.700 1617.000 ;
    RECT 1162.980 1.400 1163.820 1617.000 ;
    RECT 1164.100 1.400 1164.940 1617.000 ;
    RECT 1165.220 1.400 1166.060 1617.000 ;
    RECT 1166.340 1.400 1167.180 1617.000 ;
    RECT 1167.460 1.400 1168.300 1617.000 ;
    RECT 1168.580 1.400 1169.420 1617.000 ;
    RECT 1169.700 1.400 1170.540 1617.000 ;
    RECT 1170.820 1.400 1171.660 1617.000 ;
    RECT 1171.940 1.400 1172.780 1617.000 ;
    RECT 1173.060 1.400 1173.900 1617.000 ;
    RECT 1174.180 1.400 1175.020 1617.000 ;
    RECT 1175.300 1.400 1176.140 1617.000 ;
    RECT 1176.420 1.400 1177.260 1617.000 ;
    RECT 1177.540 1.400 1178.380 1617.000 ;
    RECT 1178.660 1.400 1179.500 1617.000 ;
    RECT 1179.780 1.400 1180.620 1617.000 ;
    RECT 1180.900 1.400 1181.740 1617.000 ;
    RECT 1182.020 1.400 1182.860 1617.000 ;
    RECT 1183.140 1.400 1183.980 1617.000 ;
    RECT 1184.260 1.400 1185.100 1617.000 ;
    RECT 1185.380 1.400 1186.220 1617.000 ;
    RECT 1186.500 1.400 1187.340 1617.000 ;
    RECT 1187.620 1.400 1188.460 1617.000 ;
    RECT 1188.740 1.400 1189.580 1617.000 ;
    RECT 1189.860 1.400 1190.700 1617.000 ;
    RECT 1190.980 1.400 1191.820 1617.000 ;
    RECT 1192.100 1.400 1192.940 1617.000 ;
    RECT 1193.220 1.400 1194.060 1617.000 ;
    RECT 1194.340 1.400 1195.180 1617.000 ;
    RECT 1195.460 1.400 1196.300 1617.000 ;
    RECT 1196.580 1.400 1197.420 1617.000 ;
    RECT 1197.700 1.400 1198.540 1617.000 ;
    RECT 1198.820 1.400 1199.660 1617.000 ;
    RECT 1199.940 1.400 1200.780 1617.000 ;
    RECT 1201.060 1.400 1201.900 1617.000 ;
    RECT 1202.180 1.400 1203.020 1617.000 ;
    RECT 1203.300 1.400 1204.140 1617.000 ;
    RECT 1204.420 1.400 1205.260 1617.000 ;
    RECT 1205.540 1.400 1206.380 1617.000 ;
    RECT 1206.660 1.400 1207.500 1617.000 ;
    RECT 1207.780 1.400 1208.620 1617.000 ;
    RECT 1208.900 1.400 1209.740 1617.000 ;
    RECT 1210.020 1.400 1210.860 1617.000 ;
    RECT 1211.140 1.400 1211.980 1617.000 ;
    RECT 1212.260 1.400 1213.100 1617.000 ;
    RECT 1213.380 1.400 1214.220 1617.000 ;
    RECT 1214.500 1.400 1215.340 1617.000 ;
    RECT 1215.620 1.400 1216.460 1617.000 ;
    RECT 1216.740 1.400 1217.580 1617.000 ;
    RECT 1217.860 1.400 1218.700 1617.000 ;
    RECT 1218.980 1.400 1219.820 1617.000 ;
    RECT 1220.100 1.400 1220.940 1617.000 ;
    RECT 1221.220 1.400 1222.060 1617.000 ;
    RECT 1222.340 1.400 1223.180 1617.000 ;
    RECT 1223.460 1.400 1224.300 1617.000 ;
    RECT 1224.580 1.400 1225.420 1617.000 ;
    RECT 1225.700 1.400 1226.540 1617.000 ;
    RECT 1226.820 1.400 1227.660 1617.000 ;
    RECT 1227.940 1.400 1228.780 1617.000 ;
    RECT 1229.060 1.400 1229.900 1617.000 ;
    RECT 1230.180 1.400 1231.020 1617.000 ;
    RECT 1231.300 1.400 1232.140 1617.000 ;
    RECT 1232.420 1.400 1233.260 1617.000 ;
    RECT 1233.540 1.400 1234.380 1617.000 ;
    RECT 1234.660 1.400 1235.500 1617.000 ;
    RECT 1235.780 1.400 1236.620 1617.000 ;
    RECT 1236.900 1.400 1237.740 1617.000 ;
    RECT 1238.020 1.400 1238.860 1617.000 ;
    RECT 1239.140 1.400 1239.980 1617.000 ;
    RECT 1240.260 1.400 1241.100 1617.000 ;
    RECT 1241.380 1.400 1242.220 1617.000 ;
    RECT 1242.500 1.400 1243.340 1617.000 ;
    RECT 1243.620 1.400 1244.460 1617.000 ;
    RECT 1244.740 1.400 1245.580 1617.000 ;
    RECT 1245.860 1.400 1246.700 1617.000 ;
    RECT 1246.980 1.400 1247.820 1617.000 ;
    RECT 1248.100 1.400 1248.940 1617.000 ;
    RECT 1249.220 1.400 1250.060 1617.000 ;
    RECT 1250.340 1.400 1251.180 1617.000 ;
    RECT 1251.460 1.400 1252.300 1617.000 ;
    RECT 1252.580 1.400 1253.420 1617.000 ;
    RECT 1253.700 1.400 1254.540 1617.000 ;
    RECT 1254.820 1.400 1255.660 1617.000 ;
    RECT 1255.940 1.400 1256.780 1617.000 ;
    RECT 1257.060 1.400 1257.900 1617.000 ;
    RECT 1258.180 1.400 1259.020 1617.000 ;
    RECT 1259.300 1.400 1260.140 1617.000 ;
    RECT 1260.420 1.400 1261.260 1617.000 ;
    RECT 1261.540 1.400 1262.380 1617.000 ;
    RECT 1262.660 1.400 1263.500 1617.000 ;
    RECT 1263.780 1.400 1264.620 1617.000 ;
    RECT 1264.900 1.400 1265.740 1617.000 ;
    RECT 1266.020 1.400 1266.860 1617.000 ;
    RECT 1267.140 1.400 1267.980 1617.000 ;
    RECT 1268.260 1.400 1269.100 1617.000 ;
    RECT 1269.380 1.400 1270.220 1617.000 ;
    RECT 1270.500 1.400 1271.340 1617.000 ;
    RECT 1271.620 1.400 1272.460 1617.000 ;
    RECT 1272.740 1.400 1273.580 1617.000 ;
    RECT 1273.860 1.400 1274.700 1617.000 ;
    RECT 1274.980 1.400 1275.820 1617.000 ;
    RECT 1276.100 1.400 1276.940 1617.000 ;
    RECT 1277.220 1.400 1278.060 1617.000 ;
    RECT 1278.340 1.400 1279.180 1617.000 ;
    RECT 1279.460 1.400 1280.300 1617.000 ;
    RECT 1280.580 1.400 1281.420 1617.000 ;
    RECT 1281.700 1.400 1282.540 1617.000 ;
    RECT 1282.820 1.400 1283.660 1617.000 ;
    RECT 1283.940 1.400 1284.780 1617.000 ;
    RECT 1285.060 1.400 1285.900 1617.000 ;
    RECT 1286.180 1.400 1287.020 1617.000 ;
    RECT 1287.300 1.400 1288.140 1617.000 ;
    RECT 1288.420 1.400 1289.260 1617.000 ;
    RECT 1289.540 1.400 1290.380 1617.000 ;
    RECT 1290.660 1.400 1291.500 1617.000 ;
    RECT 1291.780 1.400 1292.620 1617.000 ;
    RECT 1292.900 1.400 1293.740 1617.000 ;
    RECT 1294.020 1.400 1294.860 1617.000 ;
    RECT 1295.140 1.400 1295.980 1617.000 ;
    RECT 1296.260 1.400 1297.100 1617.000 ;
    RECT 1297.380 1.400 1298.220 1617.000 ;
    RECT 1298.500 1.400 1299.340 1617.000 ;
    RECT 1299.620 1.400 1300.460 1617.000 ;
    RECT 1300.740 1.400 1301.580 1617.000 ;
    RECT 1301.860 1.400 1302.700 1617.000 ;
    RECT 1302.980 1.400 1303.820 1617.000 ;
    RECT 1304.100 1.400 1304.940 1617.000 ;
    RECT 1305.220 1.400 1306.060 1617.000 ;
    RECT 1306.340 1.400 1307.180 1617.000 ;
    RECT 1307.460 1.400 1308.300 1617.000 ;
    RECT 1308.580 1.400 1309.420 1617.000 ;
    RECT 1309.700 1.400 1310.540 1617.000 ;
    RECT 1310.820 1.400 1311.660 1617.000 ;
    RECT 1311.940 1.400 1312.780 1617.000 ;
    RECT 1313.060 1.400 1313.900 1617.000 ;
    RECT 1314.180 1.400 1315.020 1617.000 ;
    RECT 1315.300 1.400 1316.140 1617.000 ;
    RECT 1316.420 1.400 1317.260 1617.000 ;
    RECT 1317.540 1.400 1318.380 1617.000 ;
    RECT 1318.660 1.400 1319.500 1617.000 ;
    RECT 1319.780 1.400 1320.620 1617.000 ;
    RECT 1320.900 1.400 1321.740 1617.000 ;
    RECT 1322.020 1.400 1322.860 1617.000 ;
    RECT 1323.140 1.400 1323.980 1617.000 ;
    RECT 1324.260 1.400 1325.100 1617.000 ;
    RECT 1325.380 1.400 1326.220 1617.000 ;
    RECT 1326.500 1.400 1327.340 1617.000 ;
    RECT 1327.620 1.400 1328.460 1617.000 ;
    RECT 1328.740 1.400 1329.580 1617.000 ;
    RECT 1329.860 1.400 1330.700 1617.000 ;
    RECT 1330.980 1.400 1331.820 1617.000 ;
    RECT 1332.100 1.400 1332.940 1617.000 ;
    RECT 1333.220 1.400 1334.060 1617.000 ;
    RECT 1334.340 1.400 1335.180 1617.000 ;
    RECT 1335.460 1.400 1336.300 1617.000 ;
    RECT 1336.580 1.400 1337.420 1617.000 ;
    RECT 1337.700 1.400 1338.540 1617.000 ;
    RECT 1338.820 1.400 1339.660 1617.000 ;
    RECT 1339.940 1.400 1340.780 1617.000 ;
    RECT 1341.060 1.400 1341.900 1617.000 ;
    RECT 1342.180 1.400 1343.020 1617.000 ;
    RECT 1343.300 1.400 1344.140 1617.000 ;
    RECT 1344.420 1.400 1345.260 1617.000 ;
    RECT 1345.540 1.400 1346.380 1617.000 ;
    RECT 1346.660 1.400 1347.500 1617.000 ;
    RECT 1347.780 1.400 1348.620 1617.000 ;
    RECT 1348.900 1.400 1349.740 1617.000 ;
    RECT 1350.020 1.400 1350.860 1617.000 ;
    RECT 1351.140 1.400 1351.980 1617.000 ;
    RECT 1352.260 1.400 1353.100 1617.000 ;
    RECT 1353.380 1.400 1354.220 1617.000 ;
    RECT 1354.500 1.400 1355.340 1617.000 ;
    RECT 1355.620 1.400 1356.460 1617.000 ;
    RECT 1356.740 1.400 1357.580 1617.000 ;
    RECT 1357.860 1.400 1358.700 1617.000 ;
    RECT 1358.980 1.400 1359.820 1617.000 ;
    RECT 1360.100 1.400 1360.940 1617.000 ;
    RECT 1361.220 1.400 1362.060 1617.000 ;
    RECT 1362.340 1.400 1363.180 1617.000 ;
    RECT 1363.460 1.400 1364.300 1617.000 ;
    RECT 1364.580 1.400 1365.420 1617.000 ;
    RECT 1365.700 1.400 1366.540 1617.000 ;
    RECT 1366.820 1.400 1367.660 1617.000 ;
    RECT 1367.940 1.400 1368.780 1617.000 ;
    RECT 1369.060 1.400 1369.900 1617.000 ;
    RECT 1370.180 1.400 1371.020 1617.000 ;
    RECT 1371.300 1.400 1372.140 1617.000 ;
    RECT 1372.420 1.400 1373.260 1617.000 ;
    RECT 1373.540 1.400 1374.380 1617.000 ;
    RECT 1374.660 1.400 1375.500 1617.000 ;
    RECT 1375.780 1.400 1376.620 1617.000 ;
    RECT 1376.900 1.400 1377.740 1617.000 ;
    RECT 1378.020 1.400 1378.860 1617.000 ;
    RECT 1379.140 1.400 1379.980 1617.000 ;
    RECT 1380.260 1.400 1381.100 1617.000 ;
    RECT 1381.380 1.400 1382.220 1617.000 ;
    RECT 1382.500 1.400 1383.340 1617.000 ;
    RECT 1383.620 1.400 1384.460 1617.000 ;
    RECT 1384.740 1.400 1385.580 1617.000 ;
    RECT 1385.860 1.400 1386.700 1617.000 ;
    RECT 1386.980 1.400 1387.820 1617.000 ;
    RECT 1388.100 1.400 1388.940 1617.000 ;
    RECT 1389.220 1.400 1390.060 1617.000 ;
    RECT 1390.340 1.400 1391.180 1617.000 ;
    RECT 1391.460 1.400 1392.300 1617.000 ;
    RECT 1392.580 1.400 1393.420 1617.000 ;
    RECT 1393.700 1.400 1394.540 1617.000 ;
    RECT 1394.820 1.400 1395.660 1617.000 ;
    RECT 1395.940 1.400 1396.780 1617.000 ;
    RECT 1397.060 1.400 1397.900 1617.000 ;
    RECT 1398.180 1.400 1399.020 1617.000 ;
    RECT 1399.300 1.400 1400.140 1617.000 ;
    RECT 1400.420 1.400 1401.260 1617.000 ;
    RECT 1401.540 1.400 1402.380 1617.000 ;
    RECT 1402.660 1.400 1403.500 1617.000 ;
    RECT 1403.780 1.400 1404.620 1617.000 ;
    RECT 1404.900 1.400 1405.740 1617.000 ;
    RECT 1406.020 1.400 1406.860 1617.000 ;
    RECT 1407.140 1.400 1407.980 1617.000 ;
    RECT 1408.260 1.400 1409.100 1617.000 ;
    RECT 1409.380 1.400 1410.220 1617.000 ;
    RECT 1410.500 1.400 1411.340 1617.000 ;
    RECT 1411.620 1.400 1412.460 1617.000 ;
    RECT 1412.740 1.400 1413.580 1617.000 ;
    RECT 1413.860 1.400 1414.700 1617.000 ;
    RECT 1414.980 1.400 1415.820 1617.000 ;
    RECT 1416.100 1.400 1416.940 1617.000 ;
    RECT 1417.220 1.400 1418.060 1617.000 ;
    RECT 1418.340 1.400 1419.180 1617.000 ;
    RECT 1419.460 1.400 1420.300 1617.000 ;
    RECT 1420.580 1.400 1421.420 1617.000 ;
    RECT 1421.700 1.400 1422.540 1617.000 ;
    RECT 1422.820 1.400 1423.660 1617.000 ;
    RECT 1423.940 1.400 1424.780 1617.000 ;
    RECT 1425.060 1.400 1425.900 1617.000 ;
    RECT 1426.180 1.400 1427.020 1617.000 ;
    RECT 1427.300 1.400 1428.140 1617.000 ;
    RECT 1428.420 1.400 1429.260 1617.000 ;
    RECT 1429.540 1.400 1430.380 1617.000 ;
    RECT 1430.660 1.400 1431.500 1617.000 ;
    RECT 1431.780 1.400 1432.620 1617.000 ;
    RECT 1432.900 1.400 1433.740 1617.000 ;
    RECT 1434.020 1.400 1434.860 1617.000 ;
    RECT 1435.140 1.400 1435.980 1617.000 ;
    RECT 1436.260 1.400 1437.100 1617.000 ;
    RECT 1437.380 1.400 1438.220 1617.000 ;
    RECT 1438.500 1.400 1439.340 1617.000 ;
    RECT 1439.620 1.400 1440.460 1617.000 ;
    RECT 1440.740 1.400 1441.580 1617.000 ;
    RECT 1441.860 1.400 1442.700 1617.000 ;
    RECT 1442.980 1.400 1443.820 1617.000 ;
    RECT 1444.100 1.400 1444.940 1617.000 ;
    RECT 1445.220 1.400 1446.060 1617.000 ;
    RECT 1446.340 1.400 1447.180 1617.000 ;
    RECT 1447.460 1.400 1448.300 1617.000 ;
    RECT 1448.580 1.400 1449.420 1617.000 ;
    RECT 1449.700 1.400 1450.540 1617.000 ;
    RECT 1450.820 1.400 1451.660 1617.000 ;
    RECT 1451.940 1.400 1452.780 1617.000 ;
    RECT 1453.060 1.400 1453.900 1617.000 ;
    RECT 1454.180 1.400 1455.020 1617.000 ;
    RECT 1455.300 1.400 1456.140 1617.000 ;
    RECT 1456.420 1.400 1457.260 1617.000 ;
    RECT 1457.540 1.400 1458.380 1617.000 ;
    RECT 1458.660 1.400 1459.500 1617.000 ;
    RECT 1459.780 1.400 1460.620 1617.000 ;
    RECT 1460.900 1.400 1461.740 1617.000 ;
    RECT 1462.020 1.400 1462.860 1617.000 ;
    RECT 1463.140 1.400 1463.980 1617.000 ;
    RECT 1464.260 1.400 1465.100 1617.000 ;
    RECT 1465.380 1.400 1466.220 1617.000 ;
    RECT 1466.500 1.400 1467.340 1617.000 ;
    RECT 1467.620 1.400 1468.460 1617.000 ;
    RECT 1468.740 1.400 1469.580 1617.000 ;
    RECT 1469.860 1.400 1470.700 1617.000 ;
    RECT 1470.980 1.400 1471.820 1617.000 ;
    RECT 1472.100 1.400 1472.940 1617.000 ;
    RECT 1473.220 1.400 1474.060 1617.000 ;
    RECT 1474.340 1.400 1475.180 1617.000 ;
    RECT 1475.460 1.400 1476.300 1617.000 ;
    RECT 1476.580 1.400 1477.420 1617.000 ;
    RECT 1477.700 1.400 1478.540 1617.000 ;
    RECT 1478.820 1.400 1479.660 1617.000 ;
    RECT 1479.940 1.400 1480.780 1617.000 ;
    RECT 1481.060 1.400 1481.900 1617.000 ;
    RECT 1482.180 1.400 1483.020 1617.000 ;
    RECT 1483.300 1.400 1484.140 1617.000 ;
    RECT 1484.420 1.400 1485.260 1617.000 ;
    RECT 1485.540 1.400 1486.380 1617.000 ;
    RECT 1486.660 1.400 1487.500 1617.000 ;
    RECT 1487.780 1.400 1488.620 1617.000 ;
    RECT 1488.900 1.400 1489.740 1617.000 ;
    RECT 1490.020 1.400 1490.860 1617.000 ;
    RECT 1491.140 1.400 1491.980 1617.000 ;
    RECT 1492.260 1.400 1493.100 1617.000 ;
    RECT 1493.380 1.400 1494.220 1617.000 ;
    RECT 1494.500 1.400 1495.340 1617.000 ;
    RECT 1495.620 1.400 1496.460 1617.000 ;
    RECT 1496.740 1.400 1497.580 1617.000 ;
    RECT 1497.860 1.400 1498.700 1617.000 ;
    RECT 1498.980 1.400 1499.820 1617.000 ;
    RECT 1500.100 1.400 1500.940 1617.000 ;
    RECT 1501.220 1.400 1502.060 1617.000 ;
    RECT 1502.340 1.400 1503.180 1617.000 ;
    RECT 1503.460 1.400 1504.300 1617.000 ;
    RECT 1504.580 1.400 1505.420 1617.000 ;
    RECT 1505.700 1.400 1506.540 1617.000 ;
    RECT 1506.820 1.400 1507.660 1617.000 ;
    RECT 1507.940 1.400 1508.780 1617.000 ;
    RECT 1509.060 1.400 1509.900 1617.000 ;
    RECT 1510.180 1.400 1511.020 1617.000 ;
    RECT 1511.300 1.400 1512.140 1617.000 ;
    RECT 1512.420 1.400 1513.260 1617.000 ;
    RECT 1513.540 1.400 1514.380 1617.000 ;
    RECT 1514.660 1.400 1515.500 1617.000 ;
    RECT 1515.780 1.400 1516.620 1617.000 ;
    RECT 1516.900 1.400 1517.740 1617.000 ;
    RECT 1518.020 1.400 1518.860 1617.000 ;
    RECT 1519.140 1.400 1519.980 1617.000 ;
    RECT 1520.260 1.400 1521.100 1617.000 ;
    RECT 1521.380 1.400 1522.220 1617.000 ;
    RECT 1522.500 1.400 1523.340 1617.000 ;
    RECT 1523.620 1.400 1524.460 1617.000 ;
    RECT 1524.740 1.400 1525.580 1617.000 ;
    RECT 1525.860 1.400 1526.700 1617.000 ;
    RECT 1526.980 1.400 1527.820 1617.000 ;
    RECT 1528.100 1.400 1528.940 1617.000 ;
    RECT 1529.220 1.400 1530.060 1617.000 ;
    RECT 1530.340 1.400 1531.180 1617.000 ;
    RECT 1531.460 1.400 1532.300 1617.000 ;
    RECT 1532.580 1.400 1533.420 1617.000 ;
    RECT 1533.700 1.400 1534.540 1617.000 ;
    RECT 1534.820 1.400 1535.660 1617.000 ;
    RECT 1535.940 1.400 1536.780 1617.000 ;
    RECT 1537.060 1.400 1537.900 1617.000 ;
    RECT 1538.180 1.400 1539.020 1617.000 ;
    RECT 1539.300 1.400 1540.140 1617.000 ;
    RECT 1540.420 1.400 1541.260 1617.000 ;
    RECT 1541.540 1.400 1542.380 1617.000 ;
    RECT 1542.660 1.400 1543.500 1617.000 ;
    RECT 1543.780 1.400 1544.620 1617.000 ;
    RECT 1544.900 1.400 1545.740 1617.000 ;
    RECT 1546.020 1.400 1546.860 1617.000 ;
    RECT 1547.140 1.400 1547.980 1617.000 ;
    RECT 1548.260 1.400 1549.100 1617.000 ;
    RECT 1549.380 1.400 1550.220 1617.000 ;
    RECT 1550.500 1.400 1551.340 1617.000 ;
    RECT 1551.620 1.400 1552.460 1617.000 ;
    RECT 1552.740 1.400 1553.580 1617.000 ;
    RECT 1553.860 1.400 1554.700 1617.000 ;
    RECT 1554.980 1.400 1555.820 1617.000 ;
    RECT 1556.100 1.400 1556.940 1617.000 ;
    RECT 1557.220 1.400 1558.060 1617.000 ;
    RECT 1558.340 1.400 1559.180 1617.000 ;
    RECT 1559.460 1.400 1560.300 1617.000 ;
    RECT 1560.580 1.400 1561.420 1617.000 ;
    RECT 1561.700 1.400 1562.540 1617.000 ;
    RECT 1562.820 1.400 1563.660 1617.000 ;
    RECT 1563.940 1.400 1564.780 1617.000 ;
    RECT 1565.060 1.400 1565.900 1617.000 ;
    RECT 1566.180 1.400 1567.020 1617.000 ;
    RECT 1567.300 1.400 1568.140 1617.000 ;
    RECT 1568.420 1.400 1569.260 1617.000 ;
    RECT 1569.540 1.400 1570.380 1617.000 ;
    RECT 1570.660 1.400 1571.500 1617.000 ;
    RECT 1571.780 1.400 1572.620 1617.000 ;
    RECT 1572.900 1.400 1573.740 1617.000 ;
    RECT 1574.020 1.400 1574.860 1617.000 ;
    RECT 1575.140 1.400 1575.980 1617.000 ;
    RECT 1576.260 1.400 1577.100 1617.000 ;
    RECT 1577.380 1.400 1578.220 1617.000 ;
    RECT 1578.500 1.400 1579.340 1617.000 ;
    RECT 1579.620 1.400 1580.460 1617.000 ;
    RECT 1580.740 1.400 1581.580 1617.000 ;
    RECT 1581.860 1.400 1582.700 1617.000 ;
    RECT 1582.980 1.400 1583.820 1617.000 ;
    RECT 1584.100 1.400 1584.940 1617.000 ;
    RECT 1585.220 1.400 1586.060 1617.000 ;
    RECT 1586.340 1.400 1587.180 1617.000 ;
    RECT 1587.460 1.400 1588.300 1617.000 ;
    RECT 1588.580 1.400 1589.420 1617.000 ;
    RECT 1589.700 1.400 1590.540 1617.000 ;
    RECT 1590.820 1.400 1591.660 1617.000 ;
    RECT 1591.940 1.400 1592.780 1617.000 ;
    RECT 1593.060 1.400 1593.900 1617.000 ;
    RECT 1594.180 1.400 1595.020 1617.000 ;
    RECT 1595.300 1.400 1596.140 1617.000 ;
    RECT 1596.420 1.400 1597.260 1617.000 ;
    RECT 1597.540 1.400 1598.380 1617.000 ;
    RECT 1598.660 1.400 1599.500 1617.000 ;
    RECT 1599.780 1.400 1600.620 1617.000 ;
    RECT 1600.900 1.400 1601.740 1617.000 ;
    RECT 1602.020 1.400 1602.860 1617.000 ;
    RECT 1603.140 1.400 1603.980 1617.000 ;
    RECT 1604.260 1.400 1605.100 1617.000 ;
    RECT 1605.380 1.400 1606.220 1617.000 ;
    RECT 1606.500 1.400 1607.340 1617.000 ;
    RECT 1607.620 1.400 1608.460 1617.000 ;
    RECT 1608.740 1.400 1609.580 1617.000 ;
    RECT 1609.860 1.400 1610.700 1617.000 ;
    RECT 1610.980 1.400 1611.820 1617.000 ;
    RECT 1612.100 1.400 1612.940 1617.000 ;
    RECT 1613.220 1.400 1614.060 1617.000 ;
    RECT 1614.340 1.400 1615.180 1617.000 ;
    RECT 1615.460 1.400 1616.300 1617.000 ;
    RECT 1616.580 1.400 1617.420 1617.000 ;
    RECT 1617.700 1.400 1618.540 1617.000 ;
    RECT 1618.820 1.400 1619.660 1617.000 ;
    RECT 1619.940 1.400 1620.780 1617.000 ;
    RECT 1621.060 1.400 1621.900 1617.000 ;
    RECT 1622.180 1.400 1623.020 1617.000 ;
    RECT 1623.300 1.400 1624.140 1617.000 ;
    RECT 1624.420 1.400 1625.260 1617.000 ;
    RECT 1625.540 1.400 1626.380 1617.000 ;
    RECT 1626.660 1.400 1627.500 1617.000 ;
    RECT 1627.780 1.400 1628.620 1617.000 ;
    RECT 1628.900 1.400 1629.740 1617.000 ;
    RECT 1630.020 1.400 1630.860 1617.000 ;
    RECT 1631.140 1.400 1631.980 1617.000 ;
    RECT 1632.260 1.400 1633.100 1617.000 ;
    RECT 1633.380 1.400 1634.220 1617.000 ;
    RECT 1634.500 1.400 1635.340 1617.000 ;
    RECT 1635.620 1.400 1636.460 1617.000 ;
    RECT 1636.740 1.400 1637.580 1617.000 ;
    RECT 1637.860 1.400 1638.700 1617.000 ;
    RECT 1638.980 1.400 1639.820 1617.000 ;
    RECT 1640.100 1.400 1640.940 1617.000 ;
    RECT 1641.220 1.400 1642.060 1617.000 ;
    RECT 1642.340 1.400 1643.180 1617.000 ;
    RECT 1643.460 1.400 1644.300 1617.000 ;
    RECT 1644.580 1.400 1645.420 1617.000 ;
    RECT 1645.700 1.400 1646.540 1617.000 ;
    RECT 1646.820 1.400 1647.660 1617.000 ;
    RECT 1647.940 1.400 1648.780 1617.000 ;
    RECT 1649.060 1.400 1649.900 1617.000 ;
    RECT 1650.180 1.400 1651.020 1617.000 ;
    RECT 1651.300 1.400 1652.140 1617.000 ;
    RECT 1652.420 1.400 1653.260 1617.000 ;
    RECT 1653.540 1.400 1654.380 1617.000 ;
    RECT 1654.660 1.400 1655.500 1617.000 ;
    RECT 1655.780 1.400 1656.620 1617.000 ;
    RECT 1656.900 1.400 1657.740 1617.000 ;
    RECT 1658.020 1.400 1658.860 1617.000 ;
    RECT 1659.140 1.400 1659.980 1617.000 ;
    RECT 1660.260 1.400 1661.100 1617.000 ;
    RECT 1661.380 1.400 1662.220 1617.000 ;
    RECT 1662.500 1.400 1663.340 1617.000 ;
    RECT 1663.620 1.400 1664.460 1617.000 ;
    RECT 1664.740 1.400 1665.580 1617.000 ;
    RECT 1665.860 1.400 1666.700 1617.000 ;
    RECT 1666.980 1.400 1667.820 1617.000 ;
    RECT 1668.100 1.400 1668.940 1617.000 ;
    RECT 1669.220 1.400 1670.060 1617.000 ;
    RECT 1670.340 1.400 1671.180 1617.000 ;
    RECT 1671.460 1.400 1672.300 1617.000 ;
    RECT 1672.580 1.400 1673.420 1617.000 ;
    RECT 1673.700 1.400 1674.540 1617.000 ;
    RECT 1674.820 1.400 1675.660 1617.000 ;
    RECT 1675.940 1.400 1676.780 1617.000 ;
    RECT 1677.060 1.400 1677.900 1617.000 ;
    RECT 1678.180 1.400 1679.020 1617.000 ;
    RECT 1679.300 1.400 1680.140 1617.000 ;
    RECT 1680.420 1.400 1681.260 1617.000 ;
    RECT 1681.540 1.400 1682.380 1617.000 ;
    RECT 1682.660 1.400 1683.500 1617.000 ;
    RECT 1683.780 1.400 1684.620 1617.000 ;
    RECT 1684.900 1.400 1685.740 1617.000 ;
    RECT 1686.020 1.400 1686.860 1617.000 ;
    RECT 1687.140 1.400 1687.980 1617.000 ;
    RECT 1688.260 1.400 1689.100 1617.000 ;
    RECT 1689.380 1.400 1690.220 1617.000 ;
    RECT 1690.500 1.400 1691.340 1617.000 ;
    RECT 1691.620 1.400 1692.460 1617.000 ;
    RECT 1692.740 1.400 1693.580 1617.000 ;
    RECT 1693.860 1.400 1694.700 1617.000 ;
    RECT 1694.980 1.400 1695.820 1617.000 ;
    RECT 1696.100 1.400 1696.940 1617.000 ;
    RECT 1697.220 1.400 1698.060 1617.000 ;
    RECT 1698.340 1.400 1699.180 1617.000 ;
    RECT 1699.460 1.400 1700.300 1617.000 ;
    RECT 1700.580 1.400 1701.420 1617.000 ;
    RECT 1701.700 1.400 1702.540 1617.000 ;
    RECT 1702.820 1.400 1703.660 1617.000 ;
    RECT 1703.940 1.400 1704.780 1617.000 ;
    RECT 1705.060 1.400 1705.900 1617.000 ;
    RECT 1706.180 1.400 1707.020 1617.000 ;
    RECT 1707.300 1.400 1708.140 1617.000 ;
    RECT 1708.420 1.400 1709.260 1617.000 ;
    RECT 1709.540 1.400 1710.380 1617.000 ;
    RECT 1710.660 1.400 1711.500 1617.000 ;
    RECT 1711.780 1.400 1712.620 1617.000 ;
    RECT 1712.900 1.400 1713.740 1617.000 ;
    RECT 1714.020 1.400 1714.860 1617.000 ;
    RECT 1715.140 1.400 1715.980 1617.000 ;
    RECT 1716.260 1.400 1717.100 1617.000 ;
    RECT 1717.380 1.400 1718.220 1617.000 ;
    RECT 1718.500 1.400 1719.340 1617.000 ;
    RECT 1719.620 1.400 1720.460 1617.000 ;
    RECT 1720.740 1.400 1721.580 1617.000 ;
    RECT 1721.860 1.400 1722.700 1617.000 ;
    RECT 1722.980 1.400 1723.820 1617.000 ;
    RECT 1724.100 1.400 1724.940 1617.000 ;
    RECT 1725.220 1.400 1726.060 1617.000 ;
    RECT 1726.340 1.400 1727.180 1617.000 ;
    RECT 1727.460 1.400 1728.300 1617.000 ;
    RECT 1728.580 1.400 1729.420 1617.000 ;
    RECT 1729.700 1.400 1730.540 1617.000 ;
    RECT 1730.820 1.400 1731.660 1617.000 ;
    RECT 1731.940 1.400 1732.780 1617.000 ;
    RECT 1733.060 1.400 1733.900 1617.000 ;
    RECT 1734.180 1.400 1735.020 1617.000 ;
    RECT 1735.300 1.400 1736.140 1617.000 ;
    RECT 1736.420 1.400 1737.260 1617.000 ;
    RECT 1737.540 1.400 1738.380 1617.000 ;
    RECT 1738.660 1.400 1739.500 1617.000 ;
    RECT 1739.780 1.400 1740.620 1617.000 ;
    RECT 1740.900 1.400 1741.740 1617.000 ;
    RECT 1742.020 1.400 1742.860 1617.000 ;
    RECT 1743.140 1.400 1743.980 1617.000 ;
    RECT 1744.260 1.400 1745.100 1617.000 ;
    RECT 1745.380 1.400 1746.220 1617.000 ;
    RECT 1746.500 1.400 1747.340 1617.000 ;
    RECT 1747.620 1.400 1748.460 1617.000 ;
    RECT 1748.740 1.400 1749.580 1617.000 ;
    RECT 1749.860 1.400 1750.700 1617.000 ;
    RECT 1750.980 1.400 1751.820 1617.000 ;
    RECT 1752.100 1.400 1752.940 1617.000 ;
    RECT 1753.220 1.400 1754.060 1617.000 ;
    RECT 1754.340 1.400 1755.180 1617.000 ;
    RECT 1755.460 1.400 1756.300 1617.000 ;
    RECT 1756.580 1.400 1757.420 1617.000 ;
    RECT 1757.700 1.400 1758.540 1617.000 ;
    RECT 1758.820 1.400 1759.660 1617.000 ;
    RECT 1759.940 1.400 1760.780 1617.000 ;
    RECT 1761.060 1.400 1761.900 1617.000 ;
    RECT 1762.180 1.400 1763.020 1617.000 ;
    RECT 1763.300 1.400 1764.140 1617.000 ;
    RECT 1764.420 1.400 1765.260 1617.000 ;
    RECT 1765.540 1.400 1766.380 1617.000 ;
    RECT 1766.660 1.400 1767.500 1617.000 ;
    RECT 1767.780 1.400 1768.620 1617.000 ;
    RECT 1768.900 1.400 1769.740 1617.000 ;
    RECT 1770.020 1.400 1770.860 1617.000 ;
    RECT 1771.140 1.400 1771.980 1617.000 ;
    RECT 1772.260 1.400 1773.100 1617.000 ;
    RECT 1773.380 1.400 1774.220 1617.000 ;
    RECT 1774.500 1.400 1775.340 1617.000 ;
    RECT 1775.620 1.400 1776.460 1617.000 ;
    RECT 1776.740 1.400 1777.580 1617.000 ;
    RECT 1777.860 1.400 1778.700 1617.000 ;
    RECT 1778.980 1.400 1779.820 1617.000 ;
    RECT 1780.100 1.400 1780.940 1617.000 ;
    RECT 1781.220 1.400 1782.060 1617.000 ;
    RECT 1782.340 1.400 1783.180 1617.000 ;
    RECT 1783.460 1.400 1784.300 1617.000 ;
    RECT 1784.580 1.400 1785.420 1617.000 ;
    RECT 1785.700 1.400 1786.540 1617.000 ;
    RECT 1786.820 1.400 1787.660 1617.000 ;
    RECT 1787.940 1.400 1788.780 1617.000 ;
    RECT 1789.060 1.400 1789.900 1617.000 ;
    RECT 1790.180 1.400 1791.020 1617.000 ;
    RECT 1791.300 1.400 1792.140 1617.000 ;
    RECT 1792.420 1.400 1793.260 1617.000 ;
    RECT 1793.540 1.400 1794.380 1617.000 ;
    RECT 1794.660 1.400 1795.500 1617.000 ;
    RECT 1795.780 1.400 1796.620 1617.000 ;
    RECT 1796.900 1.400 1797.740 1617.000 ;
    RECT 1798.020 1.400 1798.860 1617.000 ;
    RECT 1799.140 1.400 1799.980 1617.000 ;
    RECT 1800.260 1.400 1801.100 1617.000 ;
    RECT 1801.380 1.400 1802.220 1617.000 ;
    RECT 1802.500 1.400 1803.340 1617.000 ;
    RECT 1803.620 1.400 1804.460 1617.000 ;
    RECT 1804.740 1.400 1805.580 1617.000 ;
    RECT 1805.860 1.400 1806.700 1617.000 ;
    RECT 1806.980 1.400 1807.820 1617.000 ;
    RECT 1808.100 1.400 1808.940 1617.000 ;
    RECT 1809.220 1.400 1810.060 1617.000 ;
    RECT 1810.340 1.400 1811.180 1617.000 ;
    RECT 1811.460 1.400 1812.300 1617.000 ;
    RECT 1812.580 1.400 1813.420 1617.000 ;
    RECT 1813.700 1.400 1814.540 1617.000 ;
    RECT 1814.820 1.400 1815.660 1617.000 ;
    RECT 1815.940 1.400 1816.780 1617.000 ;
    RECT 1817.060 1.400 1817.900 1617.000 ;
    RECT 1818.180 1.400 1819.020 1617.000 ;
    RECT 1819.300 1.400 1820.140 1617.000 ;
    RECT 1820.420 1.400 1821.260 1617.000 ;
    RECT 1821.540 1.400 1822.380 1617.000 ;
    RECT 1822.660 1.400 1823.500 1617.000 ;
    RECT 1823.780 1.400 1824.620 1617.000 ;
    RECT 1824.900 1.400 1825.740 1617.000 ;
    RECT 1826.020 1.400 1826.860 1617.000 ;
    RECT 1827.140 1.400 1827.980 1617.000 ;
    RECT 1828.260 1.400 1829.100 1617.000 ;
    RECT 1829.380 1.400 1830.220 1617.000 ;
    RECT 1830.500 1.400 1831.340 1617.000 ;
    RECT 1831.620 1.400 1832.460 1617.000 ;
    RECT 1832.740 1.400 1833.580 1617.000 ;
    RECT 1833.860 1.400 1834.700 1617.000 ;
    RECT 1834.980 1.400 1835.820 1617.000 ;
    RECT 1836.100 1.400 1836.940 1617.000 ;
    RECT 1837.220 1.400 1838.060 1617.000 ;
    RECT 1838.340 1.400 1839.180 1617.000 ;
    RECT 1839.460 1.400 1840.300 1617.000 ;
    RECT 1840.580 1.400 1841.420 1617.000 ;
    RECT 1841.700 1.400 1842.540 1617.000 ;
    RECT 1842.820 1.400 1843.660 1617.000 ;
    RECT 1843.940 1.400 1844.780 1617.000 ;
    RECT 1845.060 1.400 1845.900 1617.000 ;
    RECT 1846.180 1.400 1847.020 1617.000 ;
    RECT 1847.300 1.400 1848.140 1617.000 ;
    RECT 1848.420 1.400 1849.260 1617.000 ;
    RECT 1849.540 1.400 1850.380 1617.000 ;
    RECT 1850.660 1.400 1851.500 1617.000 ;
    RECT 1851.780 1.400 1852.620 1617.000 ;
    RECT 1852.900 1.400 1853.740 1617.000 ;
    RECT 1854.020 1.400 1854.860 1617.000 ;
    RECT 1855.140 1.400 1855.980 1617.000 ;
    RECT 1856.260 1.400 1857.100 1617.000 ;
    RECT 1857.380 1.400 1858.220 1617.000 ;
    RECT 1858.500 1.400 1859.340 1617.000 ;
    RECT 1859.620 1.400 1860.460 1617.000 ;
    RECT 1860.740 1.400 1861.580 1617.000 ;
    RECT 1861.860 1.400 1862.700 1617.000 ;
    RECT 1862.980 1.400 1863.820 1617.000 ;
    RECT 1864.100 1.400 1864.940 1617.000 ;
    RECT 1865.220 1.400 1866.060 1617.000 ;
    RECT 1866.340 1.400 1867.180 1617.000 ;
    RECT 1867.460 1.400 1868.300 1617.000 ;
    RECT 1868.580 1.400 1869.420 1617.000 ;
    RECT 1869.700 1.400 1870.540 1617.000 ;
    RECT 1870.820 1.400 1871.660 1617.000 ;
    RECT 1871.940 1.400 1872.780 1617.000 ;
    RECT 1873.060 1.400 1873.900 1617.000 ;
    RECT 1874.180 1.400 1875.020 1617.000 ;
    RECT 1875.300 1.400 1876.140 1617.000 ;
    RECT 1876.420 1.400 1877.260 1617.000 ;
    RECT 1877.540 1.400 1878.380 1617.000 ;
    RECT 1878.660 1.400 1879.500 1617.000 ;
    RECT 1879.780 1.400 1880.620 1617.000 ;
    RECT 1880.900 1.400 1881.740 1617.000 ;
    RECT 1882.020 1.400 1882.860 1617.000 ;
    RECT 1883.140 1.400 1883.980 1617.000 ;
    RECT 1884.260 1.400 1885.100 1617.000 ;
    RECT 1885.380 1.400 1886.220 1617.000 ;
    RECT 1886.500 1.400 1887.340 1617.000 ;
    RECT 1887.620 1.400 1888.460 1617.000 ;
    RECT 1888.740 1.400 1889.580 1617.000 ;
    RECT 1889.860 1.400 1890.700 1617.000 ;
    RECT 1890.980 1.400 1891.820 1617.000 ;
    RECT 1892.100 1.400 1892.940 1617.000 ;
    RECT 1893.220 1.400 1894.060 1617.000 ;
    RECT 1894.340 1.400 1895.180 1617.000 ;
    RECT 1895.460 1.400 1896.300 1617.000 ;
    RECT 1896.580 1.400 1897.420 1617.000 ;
    RECT 1897.700 1.400 1898.540 1617.000 ;
    RECT 1898.820 1.400 1899.660 1617.000 ;
    RECT 1899.940 1.400 1900.780 1617.000 ;
    RECT 1901.060 1.400 1901.900 1617.000 ;
    RECT 1902.180 1.400 1903.020 1617.000 ;
    RECT 1903.300 1.400 1904.140 1617.000 ;
    RECT 1904.420 1.400 1905.260 1617.000 ;
    RECT 1905.540 1.400 1906.380 1617.000 ;
    RECT 1906.660 1.400 1907.500 1617.000 ;
    RECT 1907.780 1.400 1908.620 1617.000 ;
    RECT 1908.900 1.400 1909.740 1617.000 ;
    RECT 1910.020 1.400 1910.860 1617.000 ;
    RECT 1911.140 1.400 1911.980 1617.000 ;
    RECT 1912.260 1.400 1913.100 1617.000 ;
    RECT 1913.380 1.400 1914.220 1617.000 ;
    RECT 1914.500 1.400 1915.340 1617.000 ;
    RECT 1915.620 1.400 1916.460 1617.000 ;
    RECT 1916.740 1.400 1917.580 1617.000 ;
    RECT 1917.860 1.400 1918.700 1617.000 ;
    RECT 1918.980 1.400 1919.820 1617.000 ;
    RECT 1920.100 1.400 1920.940 1617.000 ;
    RECT 1921.220 1.400 1922.060 1617.000 ;
    RECT 1922.340 1.400 1923.180 1617.000 ;
    RECT 1923.460 1.400 1924.300 1617.000 ;
    RECT 1924.580 1.400 1925.420 1617.000 ;
    RECT 1925.700 1.400 1926.540 1617.000 ;
    RECT 1926.820 1.400 1927.660 1617.000 ;
    RECT 1927.940 1.400 1928.780 1617.000 ;
    RECT 1929.060 1.400 1929.900 1617.000 ;
    RECT 1930.180 1.400 1931.020 1617.000 ;
    RECT 1931.300 1.400 1932.140 1617.000 ;
    RECT 1932.420 1.400 1933.260 1617.000 ;
    RECT 1933.540 1.400 1934.380 1617.000 ;
    RECT 1934.660 1.400 1935.500 1617.000 ;
    RECT 1935.780 1.400 1936.620 1617.000 ;
    RECT 1936.900 1.400 1937.740 1617.000 ;
    RECT 1938.020 1.400 1938.860 1617.000 ;
    RECT 1939.140 1.400 1939.980 1617.000 ;
    RECT 1940.260 1.400 1941.100 1617.000 ;
    RECT 1941.380 1.400 1942.220 1617.000 ;
    RECT 1942.500 1.400 1943.340 1617.000 ;
    RECT 1943.620 1.400 1944.460 1617.000 ;
    RECT 1944.740 1.400 1945.580 1617.000 ;
    RECT 1945.860 1.400 1946.700 1617.000 ;
    RECT 1946.980 1.400 1947.820 1617.000 ;
    RECT 1948.100 1.400 1948.940 1617.000 ;
    RECT 1949.220 1.400 1950.060 1617.000 ;
    RECT 1950.340 1.400 1951.180 1617.000 ;
    RECT 1951.460 1.400 1952.300 1617.000 ;
    RECT 1952.580 1.400 1953.420 1617.000 ;
    RECT 1953.700 1.400 1954.540 1617.000 ;
    RECT 1954.820 1.400 1955.660 1617.000 ;
    RECT 1955.940 1.400 1956.780 1617.000 ;
    RECT 1957.060 1.400 1957.900 1617.000 ;
    RECT 1958.180 1.400 1959.020 1617.000 ;
    RECT 1959.300 1.400 1960.140 1617.000 ;
    RECT 1960.420 1.400 1961.260 1617.000 ;
    RECT 1961.540 1.400 1962.380 1617.000 ;
    RECT 1962.660 1.400 1963.500 1617.000 ;
    RECT 1963.780 1.400 1964.620 1617.000 ;
    RECT 1964.900 1.400 1965.740 1617.000 ;
    RECT 1966.020 1.400 1966.860 1617.000 ;
    RECT 1967.140 1.400 1967.980 1617.000 ;
    RECT 1968.260 1.400 1969.100 1617.000 ;
    RECT 1969.380 1.400 1970.220 1617.000 ;
    RECT 1970.500 1.400 1971.340 1617.000 ;
    RECT 1971.620 1.400 1972.460 1617.000 ;
    RECT 1972.740 1.400 1973.580 1617.000 ;
    RECT 1973.860 1.400 1974.700 1617.000 ;
    RECT 1974.980 1.400 1975.820 1617.000 ;
    RECT 1976.100 1.400 1976.940 1617.000 ;
    RECT 1977.220 1.400 1978.060 1617.000 ;
    RECT 1978.340 1.400 1979.180 1617.000 ;
    RECT 1979.460 1.400 1980.300 1617.000 ;
    RECT 1980.580 1.400 1981.420 1617.000 ;
    RECT 1981.700 1.400 1982.540 1617.000 ;
    RECT 1982.820 1.400 1983.660 1617.000 ;
    RECT 1983.940 1.400 1984.780 1617.000 ;
    RECT 1985.060 1.400 1985.900 1617.000 ;
    RECT 1986.180 1.400 1987.020 1617.000 ;
    RECT 1987.300 1.400 1988.140 1617.000 ;
    RECT 1988.420 1.400 1989.260 1617.000 ;
    RECT 1989.540 1.400 1990.380 1617.000 ;
    RECT 1990.660 1.400 1991.500 1617.000 ;
    RECT 1991.780 1.400 1992.620 1617.000 ;
    RECT 1992.900 1.400 1993.740 1617.000 ;
    RECT 1994.020 1.400 1994.860 1617.000 ;
    RECT 1995.140 1.400 1995.980 1617.000 ;
    RECT 1996.260 1.400 1997.100 1617.000 ;
    RECT 1997.380 1.400 1998.220 1617.000 ;
    RECT 1998.500 1.400 1999.340 1617.000 ;
    RECT 1999.620 1.400 2000.460 1617.000 ;
    RECT 2000.740 1.400 2001.580 1617.000 ;
    RECT 2001.860 1.400 2002.700 1617.000 ;
    RECT 2002.980 1.400 2003.820 1617.000 ;
    RECT 2004.100 1.400 2004.940 1617.000 ;
    RECT 2005.220 1.400 2006.060 1617.000 ;
    RECT 2006.340 1.400 2007.180 1617.000 ;
    RECT 2007.460 1.400 2008.300 1617.000 ;
    RECT 2008.580 1.400 2009.420 1617.000 ;
    RECT 2009.700 1.400 2010.540 1617.000 ;
    RECT 2010.820 1.400 2011.660 1617.000 ;
    RECT 2011.940 1.400 2012.780 1617.000 ;
    RECT 2013.060 1.400 2013.900 1617.000 ;
    RECT 2014.180 1.400 2015.020 1617.000 ;
    RECT 2015.300 1.400 2016.140 1617.000 ;
    RECT 2016.420 1.400 2017.260 1617.000 ;
    RECT 2017.540 1.400 2018.380 1617.000 ;
    RECT 2018.660 1.400 2019.500 1617.000 ;
    RECT 2019.780 1.400 2020.620 1617.000 ;
    RECT 2020.900 1.400 2021.740 1617.000 ;
    RECT 2022.020 1.400 2022.860 1617.000 ;
    RECT 2023.140 1.400 2023.980 1617.000 ;
    RECT 2024.260 1.400 2025.100 1617.000 ;
    RECT 2025.380 1.400 2026.220 1617.000 ;
    RECT 2026.500 1.400 2027.340 1617.000 ;
    RECT 2027.620 1.400 2028.460 1617.000 ;
    RECT 2028.740 1.400 2029.580 1617.000 ;
    RECT 2029.860 1.400 2030.700 1617.000 ;
    RECT 2030.980 1.400 2031.820 1617.000 ;
    RECT 2032.100 1.400 2032.940 1617.000 ;
    RECT 2033.220 1.400 2034.060 1617.000 ;
    RECT 2034.340 1.400 2035.180 1617.000 ;
    RECT 2035.460 1.400 2036.300 1617.000 ;
    RECT 2036.580 1.400 2037.420 1617.000 ;
    RECT 2037.700 1.400 2038.540 1617.000 ;
    RECT 2038.820 1.400 2039.660 1617.000 ;
    RECT 2039.940 1.400 2040.780 1617.000 ;
    RECT 2041.060 1.400 2041.900 1617.000 ;
    RECT 2042.180 1.400 2043.020 1617.000 ;
    RECT 2043.300 1.400 2044.140 1617.000 ;
    RECT 2044.420 1.400 2045.260 1617.000 ;
    RECT 2045.540 1.400 2046.380 1617.000 ;
    RECT 2046.660 1.400 2047.500 1617.000 ;
    RECT 2047.780 1.400 2048.620 1617.000 ;
    RECT 2048.900 1.400 2049.740 1617.000 ;
    RECT 2050.020 1.400 2050.860 1617.000 ;
    RECT 2051.140 1.400 2051.980 1617.000 ;
    RECT 2052.260 1.400 2053.100 1617.000 ;
    RECT 2053.380 1.400 2054.220 1617.000 ;
    RECT 2054.500 1.400 2055.340 1617.000 ;
    RECT 2055.620 1.400 2056.460 1617.000 ;
    RECT 2056.740 1.400 2057.580 1617.000 ;
    RECT 2057.860 1.400 2058.700 1617.000 ;
    RECT 2058.980 1.400 2059.820 1617.000 ;
    RECT 2060.100 1.400 2060.940 1617.000 ;
    RECT 2061.220 1.400 2062.060 1617.000 ;
    RECT 2062.340 1.400 2063.180 1617.000 ;
    RECT 2063.460 1.400 2064.300 1617.000 ;
    RECT 2064.580 1.400 2065.420 1617.000 ;
    RECT 2065.700 1.400 2066.540 1617.000 ;
    RECT 2066.820 1.400 2067.660 1617.000 ;
    RECT 2067.940 1.400 2068.780 1617.000 ;
    RECT 2069.060 1.400 2069.900 1617.000 ;
    RECT 2070.180 1.400 2071.020 1617.000 ;
    RECT 2071.300 1.400 2072.140 1617.000 ;
    RECT 2072.420 1.400 2073.260 1617.000 ;
    RECT 2073.540 1.400 2074.380 1617.000 ;
    RECT 2074.660 1.400 2075.500 1617.000 ;
    RECT 2075.780 1.400 2076.620 1617.000 ;
    RECT 2076.900 1.400 2078.600 1617.000 ;
    LAYER OVERLAP ;
    RECT 0 0 2078.600 1618.400 ;
  END
END sram_2848x32_1rw

END LIBRARY
