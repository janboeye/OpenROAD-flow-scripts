VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO sram_64x16384_1rw
  FOREIGN sram_64x16384_1rw 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1461.480 BY 637.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.345 0.070 51.415 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.225 0.070 57.295 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.105 0.070 63.175 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.985 0.070 69.055 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.865 0.070 74.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.745 0.070 80.815 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.625 0.070 86.695 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.505 0.070 92.575 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.385 0.070 98.455 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.265 0.070 104.335 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.145 0.070 110.215 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.025 0.070 116.095 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.905 0.070 121.975 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.785 0.070 127.855 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.665 0.070 133.735 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.545 0.070 139.615 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.425 0.070 145.495 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.305 0.070 151.375 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.185 0.070 157.255 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.065 0.070 163.135 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.005 0.070 166.075 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.945 0.070 169.015 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.825 0.070 174.895 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.705 0.070 180.775 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.645 0.070 183.715 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.585 0.070 186.655 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.485 0.070 191.555 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.425 0.070 194.495 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.305 0.070 200.375 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.245 0.070 203.315 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 206.185 0.070 206.255 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.125 0.070 209.195 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 212.065 0.070 212.135 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 217.945 0.070 218.015 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 220.885 0.070 220.955 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 223.825 0.070 223.895 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.705 0.070 229.775 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.645 0.070 232.715 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.585 0.070 235.655 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.525 0.070 238.595 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.465 0.070 241.535 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.405 0.070 244.475 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 247.345 0.070 247.415 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 250.285 0.070 250.355 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 253.225 0.070 253.295 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 256.165 0.070 256.235 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.105 0.070 259.175 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.045 0.070 262.115 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.985 0.070 265.055 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.925 0.070 267.995 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 270.865 0.070 270.935 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 273.805 0.070 273.875 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 276.745 0.070 276.815 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.685 0.070 279.755 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.625 0.070 282.695 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.565 0.070 285.635 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.505 0.070 288.575 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.445 0.070 291.515 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.385 0.070 294.455 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.325 0.070 297.395 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 300.265 0.070 300.335 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 303.205 0.070 303.275 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 306.145 0.070 306.215 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.085 0.070 309.155 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.025 0.070 312.095 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.965 0.070 315.035 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.905 0.070 317.975 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.845 0.070 320.915 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 323.785 0.070 323.855 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 326.725 0.070 326.795 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 329.665 0.070 329.735 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 332.605 0.070 332.675 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 335.545 0.070 335.615 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.485 0.070 338.555 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.425 0.070 341.495 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 344.365 0.070 344.435 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 347.305 0.070 347.375 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 350.245 0.070 350.315 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.185 0.070 353.255 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.125 0.070 356.195 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 359.065 0.070 359.135 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.005 0.070 362.075 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 364.945 0.070 365.015 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.885 0.070 367.955 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 370.825 0.070 370.895 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 373.765 0.070 373.835 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 376.705 0.070 376.775 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 381.605 0.070 381.675 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 384.545 0.070 384.615 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 387.485 0.070 387.555 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 390.425 0.070 390.495 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 393.365 0.070 393.435 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 396.305 0.070 396.375 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 399.245 0.070 399.315 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 402.185 0.070 402.255 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 405.125 0.070 405.195 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 408.065 0.070 408.135 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 411.005 0.070 411.075 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 413.945 0.070 414.015 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 416.885 0.070 416.955 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 419.825 0.070 419.895 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 422.765 0.070 422.835 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 425.705 0.070 425.775 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 428.645 0.070 428.715 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 431.585 0.070 431.655 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 434.525 0.070 434.595 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 437.465 0.070 437.535 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 440.405 0.070 440.475 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 443.345 0.070 443.415 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 446.285 0.070 446.355 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 449.225 0.070 449.295 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 452.165 0.070 452.235 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 455.105 0.070 455.175 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 458.045 0.070 458.115 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 460.985 0.070 461.055 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 463.925 0.070 463.995 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 466.865 0.070 466.935 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 469.805 0.070 469.875 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 472.745 0.070 472.815 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 475.685 0.070 475.755 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 478.625 0.070 478.695 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 481.565 0.070 481.635 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 484.505 0.070 484.575 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 487.445 0.070 487.515 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 490.385 0.070 490.455 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 493.325 0.070 493.395 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 496.265 0.070 496.335 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 499.205 0.070 499.275 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 502.145 0.070 502.215 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 505.085 0.070 505.155 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 508.025 0.070 508.095 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 510.965 0.070 511.035 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 513.905 0.070 513.975 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 516.845 0.070 516.915 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 519.785 0.070 519.855 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 522.725 0.070 522.795 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 525.665 0.070 525.735 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 528.605 0.070 528.675 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 531.545 0.070 531.615 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 534.485 0.070 534.555 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 537.425 0.070 537.495 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 540.365 0.070 540.435 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 543.305 0.070 543.375 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 546.245 0.070 546.315 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 549.185 0.070 549.255 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 552.125 0.070 552.195 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 555.065 0.070 555.135 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 558.005 0.070 558.075 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 560.945 0.070 561.015 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 563.885 0.070 563.955 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 566.825 0.070 566.895 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 571.725 0.070 571.795 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 574.665 0.070 574.735 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 577.605 0.070 577.675 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 580.545 0.070 580.615 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 583.485 0.070 583.555 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 586.425 0.070 586.495 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 589.365 0.070 589.435 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 592.305 0.070 592.375 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 595.245 0.070 595.315 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 598.185 0.070 598.255 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 601.125 0.070 601.195 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 604.065 0.070 604.135 ;
    END
  END addr_in[11]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 607.005 0.070 607.075 ;
    END
  END addr_in[12]
  PIN addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 609.945 0.070 610.015 ;
    END
  END addr_in[13]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 614.845 0.070 614.915 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 617.785 0.070 617.855 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 620.725 0.070 620.795 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 635.600 ;
      RECT 3.500 1.400 3.780 635.600 ;
      RECT 5.740 1.400 6.020 635.600 ;
      RECT 7.980 1.400 8.260 635.600 ;
      RECT 10.220 1.400 10.500 635.600 ;
      RECT 12.460 1.400 12.740 635.600 ;
      RECT 14.700 1.400 14.980 635.600 ;
      RECT 16.940 1.400 17.220 635.600 ;
      RECT 19.180 1.400 19.460 635.600 ;
      RECT 21.420 1.400 21.700 635.600 ;
      RECT 23.660 1.400 23.940 635.600 ;
      RECT 25.900 1.400 26.180 635.600 ;
      RECT 28.140 1.400 28.420 635.600 ;
      RECT 30.380 1.400 30.660 635.600 ;
      RECT 32.620 1.400 32.900 635.600 ;
      RECT 34.860 1.400 35.140 635.600 ;
      RECT 37.100 1.400 37.380 635.600 ;
      RECT 39.340 1.400 39.620 635.600 ;
      RECT 41.580 1.400 41.860 635.600 ;
      RECT 43.820 1.400 44.100 635.600 ;
      RECT 46.060 1.400 46.340 635.600 ;
      RECT 48.300 1.400 48.580 635.600 ;
      RECT 50.540 1.400 50.820 635.600 ;
      RECT 52.780 1.400 53.060 635.600 ;
      RECT 55.020 1.400 55.300 635.600 ;
      RECT 57.260 1.400 57.540 635.600 ;
      RECT 59.500 1.400 59.780 635.600 ;
      RECT 61.740 1.400 62.020 635.600 ;
      RECT 63.980 1.400 64.260 635.600 ;
      RECT 66.220 1.400 66.500 635.600 ;
      RECT 68.460 1.400 68.740 635.600 ;
      RECT 70.700 1.400 70.980 635.600 ;
      RECT 72.940 1.400 73.220 635.600 ;
      RECT 75.180 1.400 75.460 635.600 ;
      RECT 77.420 1.400 77.700 635.600 ;
      RECT 79.660 1.400 79.940 635.600 ;
      RECT 81.900 1.400 82.180 635.600 ;
      RECT 84.140 1.400 84.420 635.600 ;
      RECT 86.380 1.400 86.660 635.600 ;
      RECT 88.620 1.400 88.900 635.600 ;
      RECT 90.860 1.400 91.140 635.600 ;
      RECT 93.100 1.400 93.380 635.600 ;
      RECT 95.340 1.400 95.620 635.600 ;
      RECT 97.580 1.400 97.860 635.600 ;
      RECT 99.820 1.400 100.100 635.600 ;
      RECT 102.060 1.400 102.340 635.600 ;
      RECT 104.300 1.400 104.580 635.600 ;
      RECT 106.540 1.400 106.820 635.600 ;
      RECT 108.780 1.400 109.060 635.600 ;
      RECT 111.020 1.400 111.300 635.600 ;
      RECT 113.260 1.400 113.540 635.600 ;
      RECT 115.500 1.400 115.780 635.600 ;
      RECT 117.740 1.400 118.020 635.600 ;
      RECT 119.980 1.400 120.260 635.600 ;
      RECT 122.220 1.400 122.500 635.600 ;
      RECT 124.460 1.400 124.740 635.600 ;
      RECT 126.700 1.400 126.980 635.600 ;
      RECT 128.940 1.400 129.220 635.600 ;
      RECT 131.180 1.400 131.460 635.600 ;
      RECT 133.420 1.400 133.700 635.600 ;
      RECT 135.660 1.400 135.940 635.600 ;
      RECT 137.900 1.400 138.180 635.600 ;
      RECT 140.140 1.400 140.420 635.600 ;
      RECT 142.380 1.400 142.660 635.600 ;
      RECT 144.620 1.400 144.900 635.600 ;
      RECT 146.860 1.400 147.140 635.600 ;
      RECT 149.100 1.400 149.380 635.600 ;
      RECT 151.340 1.400 151.620 635.600 ;
      RECT 153.580 1.400 153.860 635.600 ;
      RECT 155.820 1.400 156.100 635.600 ;
      RECT 158.060 1.400 158.340 635.600 ;
      RECT 160.300 1.400 160.580 635.600 ;
      RECT 162.540 1.400 162.820 635.600 ;
      RECT 164.780 1.400 165.060 635.600 ;
      RECT 167.020 1.400 167.300 635.600 ;
      RECT 169.260 1.400 169.540 635.600 ;
      RECT 171.500 1.400 171.780 635.600 ;
      RECT 173.740 1.400 174.020 635.600 ;
      RECT 175.980 1.400 176.260 635.600 ;
      RECT 178.220 1.400 178.500 635.600 ;
      RECT 180.460 1.400 180.740 635.600 ;
      RECT 182.700 1.400 182.980 635.600 ;
      RECT 184.940 1.400 185.220 635.600 ;
      RECT 187.180 1.400 187.460 635.600 ;
      RECT 189.420 1.400 189.700 635.600 ;
      RECT 191.660 1.400 191.940 635.600 ;
      RECT 193.900 1.400 194.180 635.600 ;
      RECT 196.140 1.400 196.420 635.600 ;
      RECT 198.380 1.400 198.660 635.600 ;
      RECT 200.620 1.400 200.900 635.600 ;
      RECT 202.860 1.400 203.140 635.600 ;
      RECT 205.100 1.400 205.380 635.600 ;
      RECT 207.340 1.400 207.620 635.600 ;
      RECT 209.580 1.400 209.860 635.600 ;
      RECT 211.820 1.400 212.100 635.600 ;
      RECT 214.060 1.400 214.340 635.600 ;
      RECT 216.300 1.400 216.580 635.600 ;
      RECT 218.540 1.400 218.820 635.600 ;
      RECT 220.780 1.400 221.060 635.600 ;
      RECT 223.020 1.400 223.300 635.600 ;
      RECT 225.260 1.400 225.540 635.600 ;
      RECT 227.500 1.400 227.780 635.600 ;
      RECT 229.740 1.400 230.020 635.600 ;
      RECT 231.980 1.400 232.260 635.600 ;
      RECT 234.220 1.400 234.500 635.600 ;
      RECT 236.460 1.400 236.740 635.600 ;
      RECT 238.700 1.400 238.980 635.600 ;
      RECT 240.940 1.400 241.220 635.600 ;
      RECT 243.180 1.400 243.460 635.600 ;
      RECT 245.420 1.400 245.700 635.600 ;
      RECT 247.660 1.400 247.940 635.600 ;
      RECT 249.900 1.400 250.180 635.600 ;
      RECT 252.140 1.400 252.420 635.600 ;
      RECT 254.380 1.400 254.660 635.600 ;
      RECT 256.620 1.400 256.900 635.600 ;
      RECT 258.860 1.400 259.140 635.600 ;
      RECT 261.100 1.400 261.380 635.600 ;
      RECT 263.340 1.400 263.620 635.600 ;
      RECT 265.580 1.400 265.860 635.600 ;
      RECT 267.820 1.400 268.100 635.600 ;
      RECT 270.060 1.400 270.340 635.600 ;
      RECT 272.300 1.400 272.580 635.600 ;
      RECT 274.540 1.400 274.820 635.600 ;
      RECT 276.780 1.400 277.060 635.600 ;
      RECT 279.020 1.400 279.300 635.600 ;
      RECT 281.260 1.400 281.540 635.600 ;
      RECT 283.500 1.400 283.780 635.600 ;
      RECT 285.740 1.400 286.020 635.600 ;
      RECT 287.980 1.400 288.260 635.600 ;
      RECT 290.220 1.400 290.500 635.600 ;
      RECT 292.460 1.400 292.740 635.600 ;
      RECT 294.700 1.400 294.980 635.600 ;
      RECT 296.940 1.400 297.220 635.600 ;
      RECT 299.180 1.400 299.460 635.600 ;
      RECT 301.420 1.400 301.700 635.600 ;
      RECT 303.660 1.400 303.940 635.600 ;
      RECT 305.900 1.400 306.180 635.600 ;
      RECT 308.140 1.400 308.420 635.600 ;
      RECT 310.380 1.400 310.660 635.600 ;
      RECT 312.620 1.400 312.900 635.600 ;
      RECT 314.860 1.400 315.140 635.600 ;
      RECT 317.100 1.400 317.380 635.600 ;
      RECT 319.340 1.400 319.620 635.600 ;
      RECT 321.580 1.400 321.860 635.600 ;
      RECT 323.820 1.400 324.100 635.600 ;
      RECT 326.060 1.400 326.340 635.600 ;
      RECT 328.300 1.400 328.580 635.600 ;
      RECT 330.540 1.400 330.820 635.600 ;
      RECT 332.780 1.400 333.060 635.600 ;
      RECT 335.020 1.400 335.300 635.600 ;
      RECT 337.260 1.400 337.540 635.600 ;
      RECT 339.500 1.400 339.780 635.600 ;
      RECT 341.740 1.400 342.020 635.600 ;
      RECT 343.980 1.400 344.260 635.600 ;
      RECT 346.220 1.400 346.500 635.600 ;
      RECT 348.460 1.400 348.740 635.600 ;
      RECT 350.700 1.400 350.980 635.600 ;
      RECT 352.940 1.400 353.220 635.600 ;
      RECT 355.180 1.400 355.460 635.600 ;
      RECT 357.420 1.400 357.700 635.600 ;
      RECT 359.660 1.400 359.940 635.600 ;
      RECT 361.900 1.400 362.180 635.600 ;
      RECT 364.140 1.400 364.420 635.600 ;
      RECT 366.380 1.400 366.660 635.600 ;
      RECT 368.620 1.400 368.900 635.600 ;
      RECT 370.860 1.400 371.140 635.600 ;
      RECT 373.100 1.400 373.380 635.600 ;
      RECT 375.340 1.400 375.620 635.600 ;
      RECT 377.580 1.400 377.860 635.600 ;
      RECT 379.820 1.400 380.100 635.600 ;
      RECT 382.060 1.400 382.340 635.600 ;
      RECT 384.300 1.400 384.580 635.600 ;
      RECT 386.540 1.400 386.820 635.600 ;
      RECT 388.780 1.400 389.060 635.600 ;
      RECT 391.020 1.400 391.300 635.600 ;
      RECT 393.260 1.400 393.540 635.600 ;
      RECT 395.500 1.400 395.780 635.600 ;
      RECT 397.740 1.400 398.020 635.600 ;
      RECT 399.980 1.400 400.260 635.600 ;
      RECT 402.220 1.400 402.500 635.600 ;
      RECT 404.460 1.400 404.740 635.600 ;
      RECT 406.700 1.400 406.980 635.600 ;
      RECT 408.940 1.400 409.220 635.600 ;
      RECT 411.180 1.400 411.460 635.600 ;
      RECT 413.420 1.400 413.700 635.600 ;
      RECT 415.660 1.400 415.940 635.600 ;
      RECT 417.900 1.400 418.180 635.600 ;
      RECT 420.140 1.400 420.420 635.600 ;
      RECT 422.380 1.400 422.660 635.600 ;
      RECT 424.620 1.400 424.900 635.600 ;
      RECT 426.860 1.400 427.140 635.600 ;
      RECT 429.100 1.400 429.380 635.600 ;
      RECT 431.340 1.400 431.620 635.600 ;
      RECT 433.580 1.400 433.860 635.600 ;
      RECT 435.820 1.400 436.100 635.600 ;
      RECT 438.060 1.400 438.340 635.600 ;
      RECT 440.300 1.400 440.580 635.600 ;
      RECT 442.540 1.400 442.820 635.600 ;
      RECT 444.780 1.400 445.060 635.600 ;
      RECT 447.020 1.400 447.300 635.600 ;
      RECT 449.260 1.400 449.540 635.600 ;
      RECT 451.500 1.400 451.780 635.600 ;
      RECT 453.740 1.400 454.020 635.600 ;
      RECT 455.980 1.400 456.260 635.600 ;
      RECT 458.220 1.400 458.500 635.600 ;
      RECT 460.460 1.400 460.740 635.600 ;
      RECT 462.700 1.400 462.980 635.600 ;
      RECT 464.940 1.400 465.220 635.600 ;
      RECT 467.180 1.400 467.460 635.600 ;
      RECT 469.420 1.400 469.700 635.600 ;
      RECT 471.660 1.400 471.940 635.600 ;
      RECT 473.900 1.400 474.180 635.600 ;
      RECT 476.140 1.400 476.420 635.600 ;
      RECT 478.380 1.400 478.660 635.600 ;
      RECT 480.620 1.400 480.900 635.600 ;
      RECT 482.860 1.400 483.140 635.600 ;
      RECT 485.100 1.400 485.380 635.600 ;
      RECT 487.340 1.400 487.620 635.600 ;
      RECT 489.580 1.400 489.860 635.600 ;
      RECT 491.820 1.400 492.100 635.600 ;
      RECT 494.060 1.400 494.340 635.600 ;
      RECT 496.300 1.400 496.580 635.600 ;
      RECT 498.540 1.400 498.820 635.600 ;
      RECT 500.780 1.400 501.060 635.600 ;
      RECT 503.020 1.400 503.300 635.600 ;
      RECT 505.260 1.400 505.540 635.600 ;
      RECT 507.500 1.400 507.780 635.600 ;
      RECT 509.740 1.400 510.020 635.600 ;
      RECT 511.980 1.400 512.260 635.600 ;
      RECT 514.220 1.400 514.500 635.600 ;
      RECT 516.460 1.400 516.740 635.600 ;
      RECT 518.700 1.400 518.980 635.600 ;
      RECT 520.940 1.400 521.220 635.600 ;
      RECT 523.180 1.400 523.460 635.600 ;
      RECT 525.420 1.400 525.700 635.600 ;
      RECT 527.660 1.400 527.940 635.600 ;
      RECT 529.900 1.400 530.180 635.600 ;
      RECT 532.140 1.400 532.420 635.600 ;
      RECT 534.380 1.400 534.660 635.600 ;
      RECT 536.620 1.400 536.900 635.600 ;
      RECT 538.860 1.400 539.140 635.600 ;
      RECT 541.100 1.400 541.380 635.600 ;
      RECT 543.340 1.400 543.620 635.600 ;
      RECT 545.580 1.400 545.860 635.600 ;
      RECT 547.820 1.400 548.100 635.600 ;
      RECT 550.060 1.400 550.340 635.600 ;
      RECT 552.300 1.400 552.580 635.600 ;
      RECT 554.540 1.400 554.820 635.600 ;
      RECT 556.780 1.400 557.060 635.600 ;
      RECT 559.020 1.400 559.300 635.600 ;
      RECT 561.260 1.400 561.540 635.600 ;
      RECT 563.500 1.400 563.780 635.600 ;
      RECT 565.740 1.400 566.020 635.600 ;
      RECT 567.980 1.400 568.260 635.600 ;
      RECT 570.220 1.400 570.500 635.600 ;
      RECT 572.460 1.400 572.740 635.600 ;
      RECT 574.700 1.400 574.980 635.600 ;
      RECT 576.940 1.400 577.220 635.600 ;
      RECT 579.180 1.400 579.460 635.600 ;
      RECT 581.420 1.400 581.700 635.600 ;
      RECT 583.660 1.400 583.940 635.600 ;
      RECT 585.900 1.400 586.180 635.600 ;
      RECT 588.140 1.400 588.420 635.600 ;
      RECT 590.380 1.400 590.660 635.600 ;
      RECT 592.620 1.400 592.900 635.600 ;
      RECT 594.860 1.400 595.140 635.600 ;
      RECT 597.100 1.400 597.380 635.600 ;
      RECT 599.340 1.400 599.620 635.600 ;
      RECT 601.580 1.400 601.860 635.600 ;
      RECT 603.820 1.400 604.100 635.600 ;
      RECT 606.060 1.400 606.340 635.600 ;
      RECT 608.300 1.400 608.580 635.600 ;
      RECT 610.540 1.400 610.820 635.600 ;
      RECT 612.780 1.400 613.060 635.600 ;
      RECT 615.020 1.400 615.300 635.600 ;
      RECT 617.260 1.400 617.540 635.600 ;
      RECT 619.500 1.400 619.780 635.600 ;
      RECT 621.740 1.400 622.020 635.600 ;
      RECT 623.980 1.400 624.260 635.600 ;
      RECT 626.220 1.400 626.500 635.600 ;
      RECT 628.460 1.400 628.740 635.600 ;
      RECT 630.700 1.400 630.980 635.600 ;
      RECT 632.940 1.400 633.220 635.600 ;
      RECT 635.180 1.400 635.460 635.600 ;
      RECT 637.420 1.400 637.700 635.600 ;
      RECT 639.660 1.400 639.940 635.600 ;
      RECT 641.900 1.400 642.180 635.600 ;
      RECT 644.140 1.400 644.420 635.600 ;
      RECT 646.380 1.400 646.660 635.600 ;
      RECT 648.620 1.400 648.900 635.600 ;
      RECT 650.860 1.400 651.140 635.600 ;
      RECT 653.100 1.400 653.380 635.600 ;
      RECT 655.340 1.400 655.620 635.600 ;
      RECT 657.580 1.400 657.860 635.600 ;
      RECT 659.820 1.400 660.100 635.600 ;
      RECT 662.060 1.400 662.340 635.600 ;
      RECT 664.300 1.400 664.580 635.600 ;
      RECT 666.540 1.400 666.820 635.600 ;
      RECT 668.780 1.400 669.060 635.600 ;
      RECT 671.020 1.400 671.300 635.600 ;
      RECT 673.260 1.400 673.540 635.600 ;
      RECT 675.500 1.400 675.780 635.600 ;
      RECT 677.740 1.400 678.020 635.600 ;
      RECT 679.980 1.400 680.260 635.600 ;
      RECT 682.220 1.400 682.500 635.600 ;
      RECT 684.460 1.400 684.740 635.600 ;
      RECT 686.700 1.400 686.980 635.600 ;
      RECT 688.940 1.400 689.220 635.600 ;
      RECT 691.180 1.400 691.460 635.600 ;
      RECT 693.420 1.400 693.700 635.600 ;
      RECT 695.660 1.400 695.940 635.600 ;
      RECT 697.900 1.400 698.180 635.600 ;
      RECT 700.140 1.400 700.420 635.600 ;
      RECT 702.380 1.400 702.660 635.600 ;
      RECT 704.620 1.400 704.900 635.600 ;
      RECT 706.860 1.400 707.140 635.600 ;
      RECT 709.100 1.400 709.380 635.600 ;
      RECT 711.340 1.400 711.620 635.600 ;
      RECT 713.580 1.400 713.860 635.600 ;
      RECT 715.820 1.400 716.100 635.600 ;
      RECT 718.060 1.400 718.340 635.600 ;
      RECT 720.300 1.400 720.580 635.600 ;
      RECT 722.540 1.400 722.820 635.600 ;
      RECT 724.780 1.400 725.060 635.600 ;
      RECT 727.020 1.400 727.300 635.600 ;
      RECT 729.260 1.400 729.540 635.600 ;
      RECT 731.500 1.400 731.780 635.600 ;
      RECT 733.740 1.400 734.020 635.600 ;
      RECT 735.980 1.400 736.260 635.600 ;
      RECT 738.220 1.400 738.500 635.600 ;
      RECT 740.460 1.400 740.740 635.600 ;
      RECT 742.700 1.400 742.980 635.600 ;
      RECT 744.940 1.400 745.220 635.600 ;
      RECT 747.180 1.400 747.460 635.600 ;
      RECT 749.420 1.400 749.700 635.600 ;
      RECT 751.660 1.400 751.940 635.600 ;
      RECT 753.900 1.400 754.180 635.600 ;
      RECT 756.140 1.400 756.420 635.600 ;
      RECT 758.380 1.400 758.660 635.600 ;
      RECT 760.620 1.400 760.900 635.600 ;
      RECT 762.860 1.400 763.140 635.600 ;
      RECT 765.100 1.400 765.380 635.600 ;
      RECT 767.340 1.400 767.620 635.600 ;
      RECT 769.580 1.400 769.860 635.600 ;
      RECT 771.820 1.400 772.100 635.600 ;
      RECT 774.060 1.400 774.340 635.600 ;
      RECT 776.300 1.400 776.580 635.600 ;
      RECT 778.540 1.400 778.820 635.600 ;
      RECT 780.780 1.400 781.060 635.600 ;
      RECT 783.020 1.400 783.300 635.600 ;
      RECT 785.260 1.400 785.540 635.600 ;
      RECT 787.500 1.400 787.780 635.600 ;
      RECT 789.740 1.400 790.020 635.600 ;
      RECT 791.980 1.400 792.260 635.600 ;
      RECT 794.220 1.400 794.500 635.600 ;
      RECT 796.460 1.400 796.740 635.600 ;
      RECT 798.700 1.400 798.980 635.600 ;
      RECT 800.940 1.400 801.220 635.600 ;
      RECT 803.180 1.400 803.460 635.600 ;
      RECT 805.420 1.400 805.700 635.600 ;
      RECT 807.660 1.400 807.940 635.600 ;
      RECT 809.900 1.400 810.180 635.600 ;
      RECT 812.140 1.400 812.420 635.600 ;
      RECT 814.380 1.400 814.660 635.600 ;
      RECT 816.620 1.400 816.900 635.600 ;
      RECT 818.860 1.400 819.140 635.600 ;
      RECT 821.100 1.400 821.380 635.600 ;
      RECT 823.340 1.400 823.620 635.600 ;
      RECT 825.580 1.400 825.860 635.600 ;
      RECT 827.820 1.400 828.100 635.600 ;
      RECT 830.060 1.400 830.340 635.600 ;
      RECT 832.300 1.400 832.580 635.600 ;
      RECT 834.540 1.400 834.820 635.600 ;
      RECT 836.780 1.400 837.060 635.600 ;
      RECT 839.020 1.400 839.300 635.600 ;
      RECT 841.260 1.400 841.540 635.600 ;
      RECT 843.500 1.400 843.780 635.600 ;
      RECT 845.740 1.400 846.020 635.600 ;
      RECT 847.980 1.400 848.260 635.600 ;
      RECT 850.220 1.400 850.500 635.600 ;
      RECT 852.460 1.400 852.740 635.600 ;
      RECT 854.700 1.400 854.980 635.600 ;
      RECT 856.940 1.400 857.220 635.600 ;
      RECT 859.180 1.400 859.460 635.600 ;
      RECT 861.420 1.400 861.700 635.600 ;
      RECT 863.660 1.400 863.940 635.600 ;
      RECT 865.900 1.400 866.180 635.600 ;
      RECT 868.140 1.400 868.420 635.600 ;
      RECT 870.380 1.400 870.660 635.600 ;
      RECT 872.620 1.400 872.900 635.600 ;
      RECT 874.860 1.400 875.140 635.600 ;
      RECT 877.100 1.400 877.380 635.600 ;
      RECT 879.340 1.400 879.620 635.600 ;
      RECT 881.580 1.400 881.860 635.600 ;
      RECT 883.820 1.400 884.100 635.600 ;
      RECT 886.060 1.400 886.340 635.600 ;
      RECT 888.300 1.400 888.580 635.600 ;
      RECT 890.540 1.400 890.820 635.600 ;
      RECT 892.780 1.400 893.060 635.600 ;
      RECT 895.020 1.400 895.300 635.600 ;
      RECT 897.260 1.400 897.540 635.600 ;
      RECT 899.500 1.400 899.780 635.600 ;
      RECT 901.740 1.400 902.020 635.600 ;
      RECT 903.980 1.400 904.260 635.600 ;
      RECT 906.220 1.400 906.500 635.600 ;
      RECT 908.460 1.400 908.740 635.600 ;
      RECT 910.700 1.400 910.980 635.600 ;
      RECT 912.940 1.400 913.220 635.600 ;
      RECT 915.180 1.400 915.460 635.600 ;
      RECT 917.420 1.400 917.700 635.600 ;
      RECT 919.660 1.400 919.940 635.600 ;
      RECT 921.900 1.400 922.180 635.600 ;
      RECT 924.140 1.400 924.420 635.600 ;
      RECT 926.380 1.400 926.660 635.600 ;
      RECT 928.620 1.400 928.900 635.600 ;
      RECT 930.860 1.400 931.140 635.600 ;
      RECT 933.100 1.400 933.380 635.600 ;
      RECT 935.340 1.400 935.620 635.600 ;
      RECT 937.580 1.400 937.860 635.600 ;
      RECT 939.820 1.400 940.100 635.600 ;
      RECT 942.060 1.400 942.340 635.600 ;
      RECT 944.300 1.400 944.580 635.600 ;
      RECT 946.540 1.400 946.820 635.600 ;
      RECT 948.780 1.400 949.060 635.600 ;
      RECT 951.020 1.400 951.300 635.600 ;
      RECT 953.260 1.400 953.540 635.600 ;
      RECT 955.500 1.400 955.780 635.600 ;
      RECT 957.740 1.400 958.020 635.600 ;
      RECT 959.980 1.400 960.260 635.600 ;
      RECT 962.220 1.400 962.500 635.600 ;
      RECT 964.460 1.400 964.740 635.600 ;
      RECT 966.700 1.400 966.980 635.600 ;
      RECT 968.940 1.400 969.220 635.600 ;
      RECT 971.180 1.400 971.460 635.600 ;
      RECT 973.420 1.400 973.700 635.600 ;
      RECT 975.660 1.400 975.940 635.600 ;
      RECT 977.900 1.400 978.180 635.600 ;
      RECT 980.140 1.400 980.420 635.600 ;
      RECT 982.380 1.400 982.660 635.600 ;
      RECT 984.620 1.400 984.900 635.600 ;
      RECT 986.860 1.400 987.140 635.600 ;
      RECT 989.100 1.400 989.380 635.600 ;
      RECT 991.340 1.400 991.620 635.600 ;
      RECT 993.580 1.400 993.860 635.600 ;
      RECT 995.820 1.400 996.100 635.600 ;
      RECT 998.060 1.400 998.340 635.600 ;
      RECT 1000.300 1.400 1000.580 635.600 ;
      RECT 1002.540 1.400 1002.820 635.600 ;
      RECT 1004.780 1.400 1005.060 635.600 ;
      RECT 1007.020 1.400 1007.300 635.600 ;
      RECT 1009.260 1.400 1009.540 635.600 ;
      RECT 1011.500 1.400 1011.780 635.600 ;
      RECT 1013.740 1.400 1014.020 635.600 ;
      RECT 1015.980 1.400 1016.260 635.600 ;
      RECT 1018.220 1.400 1018.500 635.600 ;
      RECT 1020.460 1.400 1020.740 635.600 ;
      RECT 1022.700 1.400 1022.980 635.600 ;
      RECT 1024.940 1.400 1025.220 635.600 ;
      RECT 1027.180 1.400 1027.460 635.600 ;
      RECT 1029.420 1.400 1029.700 635.600 ;
      RECT 1031.660 1.400 1031.940 635.600 ;
      RECT 1033.900 1.400 1034.180 635.600 ;
      RECT 1036.140 1.400 1036.420 635.600 ;
      RECT 1038.380 1.400 1038.660 635.600 ;
      RECT 1040.620 1.400 1040.900 635.600 ;
      RECT 1042.860 1.400 1043.140 635.600 ;
      RECT 1045.100 1.400 1045.380 635.600 ;
      RECT 1047.340 1.400 1047.620 635.600 ;
      RECT 1049.580 1.400 1049.860 635.600 ;
      RECT 1051.820 1.400 1052.100 635.600 ;
      RECT 1054.060 1.400 1054.340 635.600 ;
      RECT 1056.300 1.400 1056.580 635.600 ;
      RECT 1058.540 1.400 1058.820 635.600 ;
      RECT 1060.780 1.400 1061.060 635.600 ;
      RECT 1063.020 1.400 1063.300 635.600 ;
      RECT 1065.260 1.400 1065.540 635.600 ;
      RECT 1067.500 1.400 1067.780 635.600 ;
      RECT 1069.740 1.400 1070.020 635.600 ;
      RECT 1071.980 1.400 1072.260 635.600 ;
      RECT 1074.220 1.400 1074.500 635.600 ;
      RECT 1076.460 1.400 1076.740 635.600 ;
      RECT 1078.700 1.400 1078.980 635.600 ;
      RECT 1080.940 1.400 1081.220 635.600 ;
      RECT 1083.180 1.400 1083.460 635.600 ;
      RECT 1085.420 1.400 1085.700 635.600 ;
      RECT 1087.660 1.400 1087.940 635.600 ;
      RECT 1089.900 1.400 1090.180 635.600 ;
      RECT 1092.140 1.400 1092.420 635.600 ;
      RECT 1094.380 1.400 1094.660 635.600 ;
      RECT 1096.620 1.400 1096.900 635.600 ;
      RECT 1098.860 1.400 1099.140 635.600 ;
      RECT 1101.100 1.400 1101.380 635.600 ;
      RECT 1103.340 1.400 1103.620 635.600 ;
      RECT 1105.580 1.400 1105.860 635.600 ;
      RECT 1107.820 1.400 1108.100 635.600 ;
      RECT 1110.060 1.400 1110.340 635.600 ;
      RECT 1112.300 1.400 1112.580 635.600 ;
      RECT 1114.540 1.400 1114.820 635.600 ;
      RECT 1116.780 1.400 1117.060 635.600 ;
      RECT 1119.020 1.400 1119.300 635.600 ;
      RECT 1121.260 1.400 1121.540 635.600 ;
      RECT 1123.500 1.400 1123.780 635.600 ;
      RECT 1125.740 1.400 1126.020 635.600 ;
      RECT 1127.980 1.400 1128.260 635.600 ;
      RECT 1130.220 1.400 1130.500 635.600 ;
      RECT 1132.460 1.400 1132.740 635.600 ;
      RECT 1134.700 1.400 1134.980 635.600 ;
      RECT 1136.940 1.400 1137.220 635.600 ;
      RECT 1139.180 1.400 1139.460 635.600 ;
      RECT 1141.420 1.400 1141.700 635.600 ;
      RECT 1143.660 1.400 1143.940 635.600 ;
      RECT 1145.900 1.400 1146.180 635.600 ;
      RECT 1148.140 1.400 1148.420 635.600 ;
      RECT 1150.380 1.400 1150.660 635.600 ;
      RECT 1152.620 1.400 1152.900 635.600 ;
      RECT 1154.860 1.400 1155.140 635.600 ;
      RECT 1157.100 1.400 1157.380 635.600 ;
      RECT 1159.340 1.400 1159.620 635.600 ;
      RECT 1161.580 1.400 1161.860 635.600 ;
      RECT 1163.820 1.400 1164.100 635.600 ;
      RECT 1166.060 1.400 1166.340 635.600 ;
      RECT 1168.300 1.400 1168.580 635.600 ;
      RECT 1170.540 1.400 1170.820 635.600 ;
      RECT 1172.780 1.400 1173.060 635.600 ;
      RECT 1175.020 1.400 1175.300 635.600 ;
      RECT 1177.260 1.400 1177.540 635.600 ;
      RECT 1179.500 1.400 1179.780 635.600 ;
      RECT 1181.740 1.400 1182.020 635.600 ;
      RECT 1183.980 1.400 1184.260 635.600 ;
      RECT 1186.220 1.400 1186.500 635.600 ;
      RECT 1188.460 1.400 1188.740 635.600 ;
      RECT 1190.700 1.400 1190.980 635.600 ;
      RECT 1192.940 1.400 1193.220 635.600 ;
      RECT 1195.180 1.400 1195.460 635.600 ;
      RECT 1197.420 1.400 1197.700 635.600 ;
      RECT 1199.660 1.400 1199.940 635.600 ;
      RECT 1201.900 1.400 1202.180 635.600 ;
      RECT 1204.140 1.400 1204.420 635.600 ;
      RECT 1206.380 1.400 1206.660 635.600 ;
      RECT 1208.620 1.400 1208.900 635.600 ;
      RECT 1210.860 1.400 1211.140 635.600 ;
      RECT 1213.100 1.400 1213.380 635.600 ;
      RECT 1215.340 1.400 1215.620 635.600 ;
      RECT 1217.580 1.400 1217.860 635.600 ;
      RECT 1219.820 1.400 1220.100 635.600 ;
      RECT 1222.060 1.400 1222.340 635.600 ;
      RECT 1224.300 1.400 1224.580 635.600 ;
      RECT 1226.540 1.400 1226.820 635.600 ;
      RECT 1228.780 1.400 1229.060 635.600 ;
      RECT 1231.020 1.400 1231.300 635.600 ;
      RECT 1233.260 1.400 1233.540 635.600 ;
      RECT 1235.500 1.400 1235.780 635.600 ;
      RECT 1237.740 1.400 1238.020 635.600 ;
      RECT 1239.980 1.400 1240.260 635.600 ;
      RECT 1242.220 1.400 1242.500 635.600 ;
      RECT 1244.460 1.400 1244.740 635.600 ;
      RECT 1246.700 1.400 1246.980 635.600 ;
      RECT 1248.940 1.400 1249.220 635.600 ;
      RECT 1251.180 1.400 1251.460 635.600 ;
      RECT 1253.420 1.400 1253.700 635.600 ;
      RECT 1255.660 1.400 1255.940 635.600 ;
      RECT 1257.900 1.400 1258.180 635.600 ;
      RECT 1260.140 1.400 1260.420 635.600 ;
      RECT 1262.380 1.400 1262.660 635.600 ;
      RECT 1264.620 1.400 1264.900 635.600 ;
      RECT 1266.860 1.400 1267.140 635.600 ;
      RECT 1269.100 1.400 1269.380 635.600 ;
      RECT 1271.340 1.400 1271.620 635.600 ;
      RECT 1273.580 1.400 1273.860 635.600 ;
      RECT 1275.820 1.400 1276.100 635.600 ;
      RECT 1278.060 1.400 1278.340 635.600 ;
      RECT 1280.300 1.400 1280.580 635.600 ;
      RECT 1282.540 1.400 1282.820 635.600 ;
      RECT 1284.780 1.400 1285.060 635.600 ;
      RECT 1287.020 1.400 1287.300 635.600 ;
      RECT 1289.260 1.400 1289.540 635.600 ;
      RECT 1291.500 1.400 1291.780 635.600 ;
      RECT 1293.740 1.400 1294.020 635.600 ;
      RECT 1295.980 1.400 1296.260 635.600 ;
      RECT 1298.220 1.400 1298.500 635.600 ;
      RECT 1300.460 1.400 1300.740 635.600 ;
      RECT 1302.700 1.400 1302.980 635.600 ;
      RECT 1304.940 1.400 1305.220 635.600 ;
      RECT 1307.180 1.400 1307.460 635.600 ;
      RECT 1309.420 1.400 1309.700 635.600 ;
      RECT 1311.660 1.400 1311.940 635.600 ;
      RECT 1313.900 1.400 1314.180 635.600 ;
      RECT 1316.140 1.400 1316.420 635.600 ;
      RECT 1318.380 1.400 1318.660 635.600 ;
      RECT 1320.620 1.400 1320.900 635.600 ;
      RECT 1322.860 1.400 1323.140 635.600 ;
      RECT 1325.100 1.400 1325.380 635.600 ;
      RECT 1327.340 1.400 1327.620 635.600 ;
      RECT 1329.580 1.400 1329.860 635.600 ;
      RECT 1331.820 1.400 1332.100 635.600 ;
      RECT 1334.060 1.400 1334.340 635.600 ;
      RECT 1336.300 1.400 1336.580 635.600 ;
      RECT 1338.540 1.400 1338.820 635.600 ;
      RECT 1340.780 1.400 1341.060 635.600 ;
      RECT 1343.020 1.400 1343.300 635.600 ;
      RECT 1345.260 1.400 1345.540 635.600 ;
      RECT 1347.500 1.400 1347.780 635.600 ;
      RECT 1349.740 1.400 1350.020 635.600 ;
      RECT 1351.980 1.400 1352.260 635.600 ;
      RECT 1354.220 1.400 1354.500 635.600 ;
      RECT 1356.460 1.400 1356.740 635.600 ;
      RECT 1358.700 1.400 1358.980 635.600 ;
      RECT 1360.940 1.400 1361.220 635.600 ;
      RECT 1363.180 1.400 1363.460 635.600 ;
      RECT 1365.420 1.400 1365.700 635.600 ;
      RECT 1367.660 1.400 1367.940 635.600 ;
      RECT 1369.900 1.400 1370.180 635.600 ;
      RECT 1372.140 1.400 1372.420 635.600 ;
      RECT 1374.380 1.400 1374.660 635.600 ;
      RECT 1376.620 1.400 1376.900 635.600 ;
      RECT 1378.860 1.400 1379.140 635.600 ;
      RECT 1381.100 1.400 1381.380 635.600 ;
      RECT 1383.340 1.400 1383.620 635.600 ;
      RECT 1385.580 1.400 1385.860 635.600 ;
      RECT 1387.820 1.400 1388.100 635.600 ;
      RECT 1390.060 1.400 1390.340 635.600 ;
      RECT 1392.300 1.400 1392.580 635.600 ;
      RECT 1394.540 1.400 1394.820 635.600 ;
      RECT 1396.780 1.400 1397.060 635.600 ;
      RECT 1399.020 1.400 1399.300 635.600 ;
      RECT 1401.260 1.400 1401.540 635.600 ;
      RECT 1403.500 1.400 1403.780 635.600 ;
      RECT 1405.740 1.400 1406.020 635.600 ;
      RECT 1407.980 1.400 1408.260 635.600 ;
      RECT 1410.220 1.400 1410.500 635.600 ;
      RECT 1412.460 1.400 1412.740 635.600 ;
      RECT 1414.700 1.400 1414.980 635.600 ;
      RECT 1416.940 1.400 1417.220 635.600 ;
      RECT 1419.180 1.400 1419.460 635.600 ;
      RECT 1421.420 1.400 1421.700 635.600 ;
      RECT 1423.660 1.400 1423.940 635.600 ;
      RECT 1425.900 1.400 1426.180 635.600 ;
      RECT 1428.140 1.400 1428.420 635.600 ;
      RECT 1430.380 1.400 1430.660 635.600 ;
      RECT 1432.620 1.400 1432.900 635.600 ;
      RECT 1434.860 1.400 1435.140 635.600 ;
      RECT 1437.100 1.400 1437.380 635.600 ;
      RECT 1439.340 1.400 1439.620 635.600 ;
      RECT 1441.580 1.400 1441.860 635.600 ;
      RECT 1443.820 1.400 1444.100 635.600 ;
      RECT 1446.060 1.400 1446.340 635.600 ;
      RECT 1448.300 1.400 1448.580 635.600 ;
      RECT 1450.540 1.400 1450.820 635.600 ;
      RECT 1452.780 1.400 1453.060 635.600 ;
      RECT 1455.020 1.400 1455.300 635.600 ;
      RECT 1457.260 1.400 1457.540 635.600 ;
      RECT 1459.500 1.400 1459.780 635.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 635.600 ;
      RECT 4.620 1.400 4.900 635.600 ;
      RECT 6.860 1.400 7.140 635.600 ;
      RECT 9.100 1.400 9.380 635.600 ;
      RECT 11.340 1.400 11.620 635.600 ;
      RECT 13.580 1.400 13.860 635.600 ;
      RECT 15.820 1.400 16.100 635.600 ;
      RECT 18.060 1.400 18.340 635.600 ;
      RECT 20.300 1.400 20.580 635.600 ;
      RECT 22.540 1.400 22.820 635.600 ;
      RECT 24.780 1.400 25.060 635.600 ;
      RECT 27.020 1.400 27.300 635.600 ;
      RECT 29.260 1.400 29.540 635.600 ;
      RECT 31.500 1.400 31.780 635.600 ;
      RECT 33.740 1.400 34.020 635.600 ;
      RECT 35.980 1.400 36.260 635.600 ;
      RECT 38.220 1.400 38.500 635.600 ;
      RECT 40.460 1.400 40.740 635.600 ;
      RECT 42.700 1.400 42.980 635.600 ;
      RECT 44.940 1.400 45.220 635.600 ;
      RECT 47.180 1.400 47.460 635.600 ;
      RECT 49.420 1.400 49.700 635.600 ;
      RECT 51.660 1.400 51.940 635.600 ;
      RECT 53.900 1.400 54.180 635.600 ;
      RECT 56.140 1.400 56.420 635.600 ;
      RECT 58.380 1.400 58.660 635.600 ;
      RECT 60.620 1.400 60.900 635.600 ;
      RECT 62.860 1.400 63.140 635.600 ;
      RECT 65.100 1.400 65.380 635.600 ;
      RECT 67.340 1.400 67.620 635.600 ;
      RECT 69.580 1.400 69.860 635.600 ;
      RECT 71.820 1.400 72.100 635.600 ;
      RECT 74.060 1.400 74.340 635.600 ;
      RECT 76.300 1.400 76.580 635.600 ;
      RECT 78.540 1.400 78.820 635.600 ;
      RECT 80.780 1.400 81.060 635.600 ;
      RECT 83.020 1.400 83.300 635.600 ;
      RECT 85.260 1.400 85.540 635.600 ;
      RECT 87.500 1.400 87.780 635.600 ;
      RECT 89.740 1.400 90.020 635.600 ;
      RECT 91.980 1.400 92.260 635.600 ;
      RECT 94.220 1.400 94.500 635.600 ;
      RECT 96.460 1.400 96.740 635.600 ;
      RECT 98.700 1.400 98.980 635.600 ;
      RECT 100.940 1.400 101.220 635.600 ;
      RECT 103.180 1.400 103.460 635.600 ;
      RECT 105.420 1.400 105.700 635.600 ;
      RECT 107.660 1.400 107.940 635.600 ;
      RECT 109.900 1.400 110.180 635.600 ;
      RECT 112.140 1.400 112.420 635.600 ;
      RECT 114.380 1.400 114.660 635.600 ;
      RECT 116.620 1.400 116.900 635.600 ;
      RECT 118.860 1.400 119.140 635.600 ;
      RECT 121.100 1.400 121.380 635.600 ;
      RECT 123.340 1.400 123.620 635.600 ;
      RECT 125.580 1.400 125.860 635.600 ;
      RECT 127.820 1.400 128.100 635.600 ;
      RECT 130.060 1.400 130.340 635.600 ;
      RECT 132.300 1.400 132.580 635.600 ;
      RECT 134.540 1.400 134.820 635.600 ;
      RECT 136.780 1.400 137.060 635.600 ;
      RECT 139.020 1.400 139.300 635.600 ;
      RECT 141.260 1.400 141.540 635.600 ;
      RECT 143.500 1.400 143.780 635.600 ;
      RECT 145.740 1.400 146.020 635.600 ;
      RECT 147.980 1.400 148.260 635.600 ;
      RECT 150.220 1.400 150.500 635.600 ;
      RECT 152.460 1.400 152.740 635.600 ;
      RECT 154.700 1.400 154.980 635.600 ;
      RECT 156.940 1.400 157.220 635.600 ;
      RECT 159.180 1.400 159.460 635.600 ;
      RECT 161.420 1.400 161.700 635.600 ;
      RECT 163.660 1.400 163.940 635.600 ;
      RECT 165.900 1.400 166.180 635.600 ;
      RECT 168.140 1.400 168.420 635.600 ;
      RECT 170.380 1.400 170.660 635.600 ;
      RECT 172.620 1.400 172.900 635.600 ;
      RECT 174.860 1.400 175.140 635.600 ;
      RECT 177.100 1.400 177.380 635.600 ;
      RECT 179.340 1.400 179.620 635.600 ;
      RECT 181.580 1.400 181.860 635.600 ;
      RECT 183.820 1.400 184.100 635.600 ;
      RECT 186.060 1.400 186.340 635.600 ;
      RECT 188.300 1.400 188.580 635.600 ;
      RECT 190.540 1.400 190.820 635.600 ;
      RECT 192.780 1.400 193.060 635.600 ;
      RECT 195.020 1.400 195.300 635.600 ;
      RECT 197.260 1.400 197.540 635.600 ;
      RECT 199.500 1.400 199.780 635.600 ;
      RECT 201.740 1.400 202.020 635.600 ;
      RECT 203.980 1.400 204.260 635.600 ;
      RECT 206.220 1.400 206.500 635.600 ;
      RECT 208.460 1.400 208.740 635.600 ;
      RECT 210.700 1.400 210.980 635.600 ;
      RECT 212.940 1.400 213.220 635.600 ;
      RECT 215.180 1.400 215.460 635.600 ;
      RECT 217.420 1.400 217.700 635.600 ;
      RECT 219.660 1.400 219.940 635.600 ;
      RECT 221.900 1.400 222.180 635.600 ;
      RECT 224.140 1.400 224.420 635.600 ;
      RECT 226.380 1.400 226.660 635.600 ;
      RECT 228.620 1.400 228.900 635.600 ;
      RECT 230.860 1.400 231.140 635.600 ;
      RECT 233.100 1.400 233.380 635.600 ;
      RECT 235.340 1.400 235.620 635.600 ;
      RECT 237.580 1.400 237.860 635.600 ;
      RECT 239.820 1.400 240.100 635.600 ;
      RECT 242.060 1.400 242.340 635.600 ;
      RECT 244.300 1.400 244.580 635.600 ;
      RECT 246.540 1.400 246.820 635.600 ;
      RECT 248.780 1.400 249.060 635.600 ;
      RECT 251.020 1.400 251.300 635.600 ;
      RECT 253.260 1.400 253.540 635.600 ;
      RECT 255.500 1.400 255.780 635.600 ;
      RECT 257.740 1.400 258.020 635.600 ;
      RECT 259.980 1.400 260.260 635.600 ;
      RECT 262.220 1.400 262.500 635.600 ;
      RECT 264.460 1.400 264.740 635.600 ;
      RECT 266.700 1.400 266.980 635.600 ;
      RECT 268.940 1.400 269.220 635.600 ;
      RECT 271.180 1.400 271.460 635.600 ;
      RECT 273.420 1.400 273.700 635.600 ;
      RECT 275.660 1.400 275.940 635.600 ;
      RECT 277.900 1.400 278.180 635.600 ;
      RECT 280.140 1.400 280.420 635.600 ;
      RECT 282.380 1.400 282.660 635.600 ;
      RECT 284.620 1.400 284.900 635.600 ;
      RECT 286.860 1.400 287.140 635.600 ;
      RECT 289.100 1.400 289.380 635.600 ;
      RECT 291.340 1.400 291.620 635.600 ;
      RECT 293.580 1.400 293.860 635.600 ;
      RECT 295.820 1.400 296.100 635.600 ;
      RECT 298.060 1.400 298.340 635.600 ;
      RECT 300.300 1.400 300.580 635.600 ;
      RECT 302.540 1.400 302.820 635.600 ;
      RECT 304.780 1.400 305.060 635.600 ;
      RECT 307.020 1.400 307.300 635.600 ;
      RECT 309.260 1.400 309.540 635.600 ;
      RECT 311.500 1.400 311.780 635.600 ;
      RECT 313.740 1.400 314.020 635.600 ;
      RECT 315.980 1.400 316.260 635.600 ;
      RECT 318.220 1.400 318.500 635.600 ;
      RECT 320.460 1.400 320.740 635.600 ;
      RECT 322.700 1.400 322.980 635.600 ;
      RECT 324.940 1.400 325.220 635.600 ;
      RECT 327.180 1.400 327.460 635.600 ;
      RECT 329.420 1.400 329.700 635.600 ;
      RECT 331.660 1.400 331.940 635.600 ;
      RECT 333.900 1.400 334.180 635.600 ;
      RECT 336.140 1.400 336.420 635.600 ;
      RECT 338.380 1.400 338.660 635.600 ;
      RECT 340.620 1.400 340.900 635.600 ;
      RECT 342.860 1.400 343.140 635.600 ;
      RECT 345.100 1.400 345.380 635.600 ;
      RECT 347.340 1.400 347.620 635.600 ;
      RECT 349.580 1.400 349.860 635.600 ;
      RECT 351.820 1.400 352.100 635.600 ;
      RECT 354.060 1.400 354.340 635.600 ;
      RECT 356.300 1.400 356.580 635.600 ;
      RECT 358.540 1.400 358.820 635.600 ;
      RECT 360.780 1.400 361.060 635.600 ;
      RECT 363.020 1.400 363.300 635.600 ;
      RECT 365.260 1.400 365.540 635.600 ;
      RECT 367.500 1.400 367.780 635.600 ;
      RECT 369.740 1.400 370.020 635.600 ;
      RECT 371.980 1.400 372.260 635.600 ;
      RECT 374.220 1.400 374.500 635.600 ;
      RECT 376.460 1.400 376.740 635.600 ;
      RECT 378.700 1.400 378.980 635.600 ;
      RECT 380.940 1.400 381.220 635.600 ;
      RECT 383.180 1.400 383.460 635.600 ;
      RECT 385.420 1.400 385.700 635.600 ;
      RECT 387.660 1.400 387.940 635.600 ;
      RECT 389.900 1.400 390.180 635.600 ;
      RECT 392.140 1.400 392.420 635.600 ;
      RECT 394.380 1.400 394.660 635.600 ;
      RECT 396.620 1.400 396.900 635.600 ;
      RECT 398.860 1.400 399.140 635.600 ;
      RECT 401.100 1.400 401.380 635.600 ;
      RECT 403.340 1.400 403.620 635.600 ;
      RECT 405.580 1.400 405.860 635.600 ;
      RECT 407.820 1.400 408.100 635.600 ;
      RECT 410.060 1.400 410.340 635.600 ;
      RECT 412.300 1.400 412.580 635.600 ;
      RECT 414.540 1.400 414.820 635.600 ;
      RECT 416.780 1.400 417.060 635.600 ;
      RECT 419.020 1.400 419.300 635.600 ;
      RECT 421.260 1.400 421.540 635.600 ;
      RECT 423.500 1.400 423.780 635.600 ;
      RECT 425.740 1.400 426.020 635.600 ;
      RECT 427.980 1.400 428.260 635.600 ;
      RECT 430.220 1.400 430.500 635.600 ;
      RECT 432.460 1.400 432.740 635.600 ;
      RECT 434.700 1.400 434.980 635.600 ;
      RECT 436.940 1.400 437.220 635.600 ;
      RECT 439.180 1.400 439.460 635.600 ;
      RECT 441.420 1.400 441.700 635.600 ;
      RECT 443.660 1.400 443.940 635.600 ;
      RECT 445.900 1.400 446.180 635.600 ;
      RECT 448.140 1.400 448.420 635.600 ;
      RECT 450.380 1.400 450.660 635.600 ;
      RECT 452.620 1.400 452.900 635.600 ;
      RECT 454.860 1.400 455.140 635.600 ;
      RECT 457.100 1.400 457.380 635.600 ;
      RECT 459.340 1.400 459.620 635.600 ;
      RECT 461.580 1.400 461.860 635.600 ;
      RECT 463.820 1.400 464.100 635.600 ;
      RECT 466.060 1.400 466.340 635.600 ;
      RECT 468.300 1.400 468.580 635.600 ;
      RECT 470.540 1.400 470.820 635.600 ;
      RECT 472.780 1.400 473.060 635.600 ;
      RECT 475.020 1.400 475.300 635.600 ;
      RECT 477.260 1.400 477.540 635.600 ;
      RECT 479.500 1.400 479.780 635.600 ;
      RECT 481.740 1.400 482.020 635.600 ;
      RECT 483.980 1.400 484.260 635.600 ;
      RECT 486.220 1.400 486.500 635.600 ;
      RECT 488.460 1.400 488.740 635.600 ;
      RECT 490.700 1.400 490.980 635.600 ;
      RECT 492.940 1.400 493.220 635.600 ;
      RECT 495.180 1.400 495.460 635.600 ;
      RECT 497.420 1.400 497.700 635.600 ;
      RECT 499.660 1.400 499.940 635.600 ;
      RECT 501.900 1.400 502.180 635.600 ;
      RECT 504.140 1.400 504.420 635.600 ;
      RECT 506.380 1.400 506.660 635.600 ;
      RECT 508.620 1.400 508.900 635.600 ;
      RECT 510.860 1.400 511.140 635.600 ;
      RECT 513.100 1.400 513.380 635.600 ;
      RECT 515.340 1.400 515.620 635.600 ;
      RECT 517.580 1.400 517.860 635.600 ;
      RECT 519.820 1.400 520.100 635.600 ;
      RECT 522.060 1.400 522.340 635.600 ;
      RECT 524.300 1.400 524.580 635.600 ;
      RECT 526.540 1.400 526.820 635.600 ;
      RECT 528.780 1.400 529.060 635.600 ;
      RECT 531.020 1.400 531.300 635.600 ;
      RECT 533.260 1.400 533.540 635.600 ;
      RECT 535.500 1.400 535.780 635.600 ;
      RECT 537.740 1.400 538.020 635.600 ;
      RECT 539.980 1.400 540.260 635.600 ;
      RECT 542.220 1.400 542.500 635.600 ;
      RECT 544.460 1.400 544.740 635.600 ;
      RECT 546.700 1.400 546.980 635.600 ;
      RECT 548.940 1.400 549.220 635.600 ;
      RECT 551.180 1.400 551.460 635.600 ;
      RECT 553.420 1.400 553.700 635.600 ;
      RECT 555.660 1.400 555.940 635.600 ;
      RECT 557.900 1.400 558.180 635.600 ;
      RECT 560.140 1.400 560.420 635.600 ;
      RECT 562.380 1.400 562.660 635.600 ;
      RECT 564.620 1.400 564.900 635.600 ;
      RECT 566.860 1.400 567.140 635.600 ;
      RECT 569.100 1.400 569.380 635.600 ;
      RECT 571.340 1.400 571.620 635.600 ;
      RECT 573.580 1.400 573.860 635.600 ;
      RECT 575.820 1.400 576.100 635.600 ;
      RECT 578.060 1.400 578.340 635.600 ;
      RECT 580.300 1.400 580.580 635.600 ;
      RECT 582.540 1.400 582.820 635.600 ;
      RECT 584.780 1.400 585.060 635.600 ;
      RECT 587.020 1.400 587.300 635.600 ;
      RECT 589.260 1.400 589.540 635.600 ;
      RECT 591.500 1.400 591.780 635.600 ;
      RECT 593.740 1.400 594.020 635.600 ;
      RECT 595.980 1.400 596.260 635.600 ;
      RECT 598.220 1.400 598.500 635.600 ;
      RECT 600.460 1.400 600.740 635.600 ;
      RECT 602.700 1.400 602.980 635.600 ;
      RECT 604.940 1.400 605.220 635.600 ;
      RECT 607.180 1.400 607.460 635.600 ;
      RECT 609.420 1.400 609.700 635.600 ;
      RECT 611.660 1.400 611.940 635.600 ;
      RECT 613.900 1.400 614.180 635.600 ;
      RECT 616.140 1.400 616.420 635.600 ;
      RECT 618.380 1.400 618.660 635.600 ;
      RECT 620.620 1.400 620.900 635.600 ;
      RECT 622.860 1.400 623.140 635.600 ;
      RECT 625.100 1.400 625.380 635.600 ;
      RECT 627.340 1.400 627.620 635.600 ;
      RECT 629.580 1.400 629.860 635.600 ;
      RECT 631.820 1.400 632.100 635.600 ;
      RECT 634.060 1.400 634.340 635.600 ;
      RECT 636.300 1.400 636.580 635.600 ;
      RECT 638.540 1.400 638.820 635.600 ;
      RECT 640.780 1.400 641.060 635.600 ;
      RECT 643.020 1.400 643.300 635.600 ;
      RECT 645.260 1.400 645.540 635.600 ;
      RECT 647.500 1.400 647.780 635.600 ;
      RECT 649.740 1.400 650.020 635.600 ;
      RECT 651.980 1.400 652.260 635.600 ;
      RECT 654.220 1.400 654.500 635.600 ;
      RECT 656.460 1.400 656.740 635.600 ;
      RECT 658.700 1.400 658.980 635.600 ;
      RECT 660.940 1.400 661.220 635.600 ;
      RECT 663.180 1.400 663.460 635.600 ;
      RECT 665.420 1.400 665.700 635.600 ;
      RECT 667.660 1.400 667.940 635.600 ;
      RECT 669.900 1.400 670.180 635.600 ;
      RECT 672.140 1.400 672.420 635.600 ;
      RECT 674.380 1.400 674.660 635.600 ;
      RECT 676.620 1.400 676.900 635.600 ;
      RECT 678.860 1.400 679.140 635.600 ;
      RECT 681.100 1.400 681.380 635.600 ;
      RECT 683.340 1.400 683.620 635.600 ;
      RECT 685.580 1.400 685.860 635.600 ;
      RECT 687.820 1.400 688.100 635.600 ;
      RECT 690.060 1.400 690.340 635.600 ;
      RECT 692.300 1.400 692.580 635.600 ;
      RECT 694.540 1.400 694.820 635.600 ;
      RECT 696.780 1.400 697.060 635.600 ;
      RECT 699.020 1.400 699.300 635.600 ;
      RECT 701.260 1.400 701.540 635.600 ;
      RECT 703.500 1.400 703.780 635.600 ;
      RECT 705.740 1.400 706.020 635.600 ;
      RECT 707.980 1.400 708.260 635.600 ;
      RECT 710.220 1.400 710.500 635.600 ;
      RECT 712.460 1.400 712.740 635.600 ;
      RECT 714.700 1.400 714.980 635.600 ;
      RECT 716.940 1.400 717.220 635.600 ;
      RECT 719.180 1.400 719.460 635.600 ;
      RECT 721.420 1.400 721.700 635.600 ;
      RECT 723.660 1.400 723.940 635.600 ;
      RECT 725.900 1.400 726.180 635.600 ;
      RECT 728.140 1.400 728.420 635.600 ;
      RECT 730.380 1.400 730.660 635.600 ;
      RECT 732.620 1.400 732.900 635.600 ;
      RECT 734.860 1.400 735.140 635.600 ;
      RECT 737.100 1.400 737.380 635.600 ;
      RECT 739.340 1.400 739.620 635.600 ;
      RECT 741.580 1.400 741.860 635.600 ;
      RECT 743.820 1.400 744.100 635.600 ;
      RECT 746.060 1.400 746.340 635.600 ;
      RECT 748.300 1.400 748.580 635.600 ;
      RECT 750.540 1.400 750.820 635.600 ;
      RECT 752.780 1.400 753.060 635.600 ;
      RECT 755.020 1.400 755.300 635.600 ;
      RECT 757.260 1.400 757.540 635.600 ;
      RECT 759.500 1.400 759.780 635.600 ;
      RECT 761.740 1.400 762.020 635.600 ;
      RECT 763.980 1.400 764.260 635.600 ;
      RECT 766.220 1.400 766.500 635.600 ;
      RECT 768.460 1.400 768.740 635.600 ;
      RECT 770.700 1.400 770.980 635.600 ;
      RECT 772.940 1.400 773.220 635.600 ;
      RECT 775.180 1.400 775.460 635.600 ;
      RECT 777.420 1.400 777.700 635.600 ;
      RECT 779.660 1.400 779.940 635.600 ;
      RECT 781.900 1.400 782.180 635.600 ;
      RECT 784.140 1.400 784.420 635.600 ;
      RECT 786.380 1.400 786.660 635.600 ;
      RECT 788.620 1.400 788.900 635.600 ;
      RECT 790.860 1.400 791.140 635.600 ;
      RECT 793.100 1.400 793.380 635.600 ;
      RECT 795.340 1.400 795.620 635.600 ;
      RECT 797.580 1.400 797.860 635.600 ;
      RECT 799.820 1.400 800.100 635.600 ;
      RECT 802.060 1.400 802.340 635.600 ;
      RECT 804.300 1.400 804.580 635.600 ;
      RECT 806.540 1.400 806.820 635.600 ;
      RECT 808.780 1.400 809.060 635.600 ;
      RECT 811.020 1.400 811.300 635.600 ;
      RECT 813.260 1.400 813.540 635.600 ;
      RECT 815.500 1.400 815.780 635.600 ;
      RECT 817.740 1.400 818.020 635.600 ;
      RECT 819.980 1.400 820.260 635.600 ;
      RECT 822.220 1.400 822.500 635.600 ;
      RECT 824.460 1.400 824.740 635.600 ;
      RECT 826.700 1.400 826.980 635.600 ;
      RECT 828.940 1.400 829.220 635.600 ;
      RECT 831.180 1.400 831.460 635.600 ;
      RECT 833.420 1.400 833.700 635.600 ;
      RECT 835.660 1.400 835.940 635.600 ;
      RECT 837.900 1.400 838.180 635.600 ;
      RECT 840.140 1.400 840.420 635.600 ;
      RECT 842.380 1.400 842.660 635.600 ;
      RECT 844.620 1.400 844.900 635.600 ;
      RECT 846.860 1.400 847.140 635.600 ;
      RECT 849.100 1.400 849.380 635.600 ;
      RECT 851.340 1.400 851.620 635.600 ;
      RECT 853.580 1.400 853.860 635.600 ;
      RECT 855.820 1.400 856.100 635.600 ;
      RECT 858.060 1.400 858.340 635.600 ;
      RECT 860.300 1.400 860.580 635.600 ;
      RECT 862.540 1.400 862.820 635.600 ;
      RECT 864.780 1.400 865.060 635.600 ;
      RECT 867.020 1.400 867.300 635.600 ;
      RECT 869.260 1.400 869.540 635.600 ;
      RECT 871.500 1.400 871.780 635.600 ;
      RECT 873.740 1.400 874.020 635.600 ;
      RECT 875.980 1.400 876.260 635.600 ;
      RECT 878.220 1.400 878.500 635.600 ;
      RECT 880.460 1.400 880.740 635.600 ;
      RECT 882.700 1.400 882.980 635.600 ;
      RECT 884.940 1.400 885.220 635.600 ;
      RECT 887.180 1.400 887.460 635.600 ;
      RECT 889.420 1.400 889.700 635.600 ;
      RECT 891.660 1.400 891.940 635.600 ;
      RECT 893.900 1.400 894.180 635.600 ;
      RECT 896.140 1.400 896.420 635.600 ;
      RECT 898.380 1.400 898.660 635.600 ;
      RECT 900.620 1.400 900.900 635.600 ;
      RECT 902.860 1.400 903.140 635.600 ;
      RECT 905.100 1.400 905.380 635.600 ;
      RECT 907.340 1.400 907.620 635.600 ;
      RECT 909.580 1.400 909.860 635.600 ;
      RECT 911.820 1.400 912.100 635.600 ;
      RECT 914.060 1.400 914.340 635.600 ;
      RECT 916.300 1.400 916.580 635.600 ;
      RECT 918.540 1.400 918.820 635.600 ;
      RECT 920.780 1.400 921.060 635.600 ;
      RECT 923.020 1.400 923.300 635.600 ;
      RECT 925.260 1.400 925.540 635.600 ;
      RECT 927.500 1.400 927.780 635.600 ;
      RECT 929.740 1.400 930.020 635.600 ;
      RECT 931.980 1.400 932.260 635.600 ;
      RECT 934.220 1.400 934.500 635.600 ;
      RECT 936.460 1.400 936.740 635.600 ;
      RECT 938.700 1.400 938.980 635.600 ;
      RECT 940.940 1.400 941.220 635.600 ;
      RECT 943.180 1.400 943.460 635.600 ;
      RECT 945.420 1.400 945.700 635.600 ;
      RECT 947.660 1.400 947.940 635.600 ;
      RECT 949.900 1.400 950.180 635.600 ;
      RECT 952.140 1.400 952.420 635.600 ;
      RECT 954.380 1.400 954.660 635.600 ;
      RECT 956.620 1.400 956.900 635.600 ;
      RECT 958.860 1.400 959.140 635.600 ;
      RECT 961.100 1.400 961.380 635.600 ;
      RECT 963.340 1.400 963.620 635.600 ;
      RECT 965.580 1.400 965.860 635.600 ;
      RECT 967.820 1.400 968.100 635.600 ;
      RECT 970.060 1.400 970.340 635.600 ;
      RECT 972.300 1.400 972.580 635.600 ;
      RECT 974.540 1.400 974.820 635.600 ;
      RECT 976.780 1.400 977.060 635.600 ;
      RECT 979.020 1.400 979.300 635.600 ;
      RECT 981.260 1.400 981.540 635.600 ;
      RECT 983.500 1.400 983.780 635.600 ;
      RECT 985.740 1.400 986.020 635.600 ;
      RECT 987.980 1.400 988.260 635.600 ;
      RECT 990.220 1.400 990.500 635.600 ;
      RECT 992.460 1.400 992.740 635.600 ;
      RECT 994.700 1.400 994.980 635.600 ;
      RECT 996.940 1.400 997.220 635.600 ;
      RECT 999.180 1.400 999.460 635.600 ;
      RECT 1001.420 1.400 1001.700 635.600 ;
      RECT 1003.660 1.400 1003.940 635.600 ;
      RECT 1005.900 1.400 1006.180 635.600 ;
      RECT 1008.140 1.400 1008.420 635.600 ;
      RECT 1010.380 1.400 1010.660 635.600 ;
      RECT 1012.620 1.400 1012.900 635.600 ;
      RECT 1014.860 1.400 1015.140 635.600 ;
      RECT 1017.100 1.400 1017.380 635.600 ;
      RECT 1019.340 1.400 1019.620 635.600 ;
      RECT 1021.580 1.400 1021.860 635.600 ;
      RECT 1023.820 1.400 1024.100 635.600 ;
      RECT 1026.060 1.400 1026.340 635.600 ;
      RECT 1028.300 1.400 1028.580 635.600 ;
      RECT 1030.540 1.400 1030.820 635.600 ;
      RECT 1032.780 1.400 1033.060 635.600 ;
      RECT 1035.020 1.400 1035.300 635.600 ;
      RECT 1037.260 1.400 1037.540 635.600 ;
      RECT 1039.500 1.400 1039.780 635.600 ;
      RECT 1041.740 1.400 1042.020 635.600 ;
      RECT 1043.980 1.400 1044.260 635.600 ;
      RECT 1046.220 1.400 1046.500 635.600 ;
      RECT 1048.460 1.400 1048.740 635.600 ;
      RECT 1050.700 1.400 1050.980 635.600 ;
      RECT 1052.940 1.400 1053.220 635.600 ;
      RECT 1055.180 1.400 1055.460 635.600 ;
      RECT 1057.420 1.400 1057.700 635.600 ;
      RECT 1059.660 1.400 1059.940 635.600 ;
      RECT 1061.900 1.400 1062.180 635.600 ;
      RECT 1064.140 1.400 1064.420 635.600 ;
      RECT 1066.380 1.400 1066.660 635.600 ;
      RECT 1068.620 1.400 1068.900 635.600 ;
      RECT 1070.860 1.400 1071.140 635.600 ;
      RECT 1073.100 1.400 1073.380 635.600 ;
      RECT 1075.340 1.400 1075.620 635.600 ;
      RECT 1077.580 1.400 1077.860 635.600 ;
      RECT 1079.820 1.400 1080.100 635.600 ;
      RECT 1082.060 1.400 1082.340 635.600 ;
      RECT 1084.300 1.400 1084.580 635.600 ;
      RECT 1086.540 1.400 1086.820 635.600 ;
      RECT 1088.780 1.400 1089.060 635.600 ;
      RECT 1091.020 1.400 1091.300 635.600 ;
      RECT 1093.260 1.400 1093.540 635.600 ;
      RECT 1095.500 1.400 1095.780 635.600 ;
      RECT 1097.740 1.400 1098.020 635.600 ;
      RECT 1099.980 1.400 1100.260 635.600 ;
      RECT 1102.220 1.400 1102.500 635.600 ;
      RECT 1104.460 1.400 1104.740 635.600 ;
      RECT 1106.700 1.400 1106.980 635.600 ;
      RECT 1108.940 1.400 1109.220 635.600 ;
      RECT 1111.180 1.400 1111.460 635.600 ;
      RECT 1113.420 1.400 1113.700 635.600 ;
      RECT 1115.660 1.400 1115.940 635.600 ;
      RECT 1117.900 1.400 1118.180 635.600 ;
      RECT 1120.140 1.400 1120.420 635.600 ;
      RECT 1122.380 1.400 1122.660 635.600 ;
      RECT 1124.620 1.400 1124.900 635.600 ;
      RECT 1126.860 1.400 1127.140 635.600 ;
      RECT 1129.100 1.400 1129.380 635.600 ;
      RECT 1131.340 1.400 1131.620 635.600 ;
      RECT 1133.580 1.400 1133.860 635.600 ;
      RECT 1135.820 1.400 1136.100 635.600 ;
      RECT 1138.060 1.400 1138.340 635.600 ;
      RECT 1140.300 1.400 1140.580 635.600 ;
      RECT 1142.540 1.400 1142.820 635.600 ;
      RECT 1144.780 1.400 1145.060 635.600 ;
      RECT 1147.020 1.400 1147.300 635.600 ;
      RECT 1149.260 1.400 1149.540 635.600 ;
      RECT 1151.500 1.400 1151.780 635.600 ;
      RECT 1153.740 1.400 1154.020 635.600 ;
      RECT 1155.980 1.400 1156.260 635.600 ;
      RECT 1158.220 1.400 1158.500 635.600 ;
      RECT 1160.460 1.400 1160.740 635.600 ;
      RECT 1162.700 1.400 1162.980 635.600 ;
      RECT 1164.940 1.400 1165.220 635.600 ;
      RECT 1167.180 1.400 1167.460 635.600 ;
      RECT 1169.420 1.400 1169.700 635.600 ;
      RECT 1171.660 1.400 1171.940 635.600 ;
      RECT 1173.900 1.400 1174.180 635.600 ;
      RECT 1176.140 1.400 1176.420 635.600 ;
      RECT 1178.380 1.400 1178.660 635.600 ;
      RECT 1180.620 1.400 1180.900 635.600 ;
      RECT 1182.860 1.400 1183.140 635.600 ;
      RECT 1185.100 1.400 1185.380 635.600 ;
      RECT 1187.340 1.400 1187.620 635.600 ;
      RECT 1189.580 1.400 1189.860 635.600 ;
      RECT 1191.820 1.400 1192.100 635.600 ;
      RECT 1194.060 1.400 1194.340 635.600 ;
      RECT 1196.300 1.400 1196.580 635.600 ;
      RECT 1198.540 1.400 1198.820 635.600 ;
      RECT 1200.780 1.400 1201.060 635.600 ;
      RECT 1203.020 1.400 1203.300 635.600 ;
      RECT 1205.260 1.400 1205.540 635.600 ;
      RECT 1207.500 1.400 1207.780 635.600 ;
      RECT 1209.740 1.400 1210.020 635.600 ;
      RECT 1211.980 1.400 1212.260 635.600 ;
      RECT 1214.220 1.400 1214.500 635.600 ;
      RECT 1216.460 1.400 1216.740 635.600 ;
      RECT 1218.700 1.400 1218.980 635.600 ;
      RECT 1220.940 1.400 1221.220 635.600 ;
      RECT 1223.180 1.400 1223.460 635.600 ;
      RECT 1225.420 1.400 1225.700 635.600 ;
      RECT 1227.660 1.400 1227.940 635.600 ;
      RECT 1229.900 1.400 1230.180 635.600 ;
      RECT 1232.140 1.400 1232.420 635.600 ;
      RECT 1234.380 1.400 1234.660 635.600 ;
      RECT 1236.620 1.400 1236.900 635.600 ;
      RECT 1238.860 1.400 1239.140 635.600 ;
      RECT 1241.100 1.400 1241.380 635.600 ;
      RECT 1243.340 1.400 1243.620 635.600 ;
      RECT 1245.580 1.400 1245.860 635.600 ;
      RECT 1247.820 1.400 1248.100 635.600 ;
      RECT 1250.060 1.400 1250.340 635.600 ;
      RECT 1252.300 1.400 1252.580 635.600 ;
      RECT 1254.540 1.400 1254.820 635.600 ;
      RECT 1256.780 1.400 1257.060 635.600 ;
      RECT 1259.020 1.400 1259.300 635.600 ;
      RECT 1261.260 1.400 1261.540 635.600 ;
      RECT 1263.500 1.400 1263.780 635.600 ;
      RECT 1265.740 1.400 1266.020 635.600 ;
      RECT 1267.980 1.400 1268.260 635.600 ;
      RECT 1270.220 1.400 1270.500 635.600 ;
      RECT 1272.460 1.400 1272.740 635.600 ;
      RECT 1274.700 1.400 1274.980 635.600 ;
      RECT 1276.940 1.400 1277.220 635.600 ;
      RECT 1279.180 1.400 1279.460 635.600 ;
      RECT 1281.420 1.400 1281.700 635.600 ;
      RECT 1283.660 1.400 1283.940 635.600 ;
      RECT 1285.900 1.400 1286.180 635.600 ;
      RECT 1288.140 1.400 1288.420 635.600 ;
      RECT 1290.380 1.400 1290.660 635.600 ;
      RECT 1292.620 1.400 1292.900 635.600 ;
      RECT 1294.860 1.400 1295.140 635.600 ;
      RECT 1297.100 1.400 1297.380 635.600 ;
      RECT 1299.340 1.400 1299.620 635.600 ;
      RECT 1301.580 1.400 1301.860 635.600 ;
      RECT 1303.820 1.400 1304.100 635.600 ;
      RECT 1306.060 1.400 1306.340 635.600 ;
      RECT 1308.300 1.400 1308.580 635.600 ;
      RECT 1310.540 1.400 1310.820 635.600 ;
      RECT 1312.780 1.400 1313.060 635.600 ;
      RECT 1315.020 1.400 1315.300 635.600 ;
      RECT 1317.260 1.400 1317.540 635.600 ;
      RECT 1319.500 1.400 1319.780 635.600 ;
      RECT 1321.740 1.400 1322.020 635.600 ;
      RECT 1323.980 1.400 1324.260 635.600 ;
      RECT 1326.220 1.400 1326.500 635.600 ;
      RECT 1328.460 1.400 1328.740 635.600 ;
      RECT 1330.700 1.400 1330.980 635.600 ;
      RECT 1332.940 1.400 1333.220 635.600 ;
      RECT 1335.180 1.400 1335.460 635.600 ;
      RECT 1337.420 1.400 1337.700 635.600 ;
      RECT 1339.660 1.400 1339.940 635.600 ;
      RECT 1341.900 1.400 1342.180 635.600 ;
      RECT 1344.140 1.400 1344.420 635.600 ;
      RECT 1346.380 1.400 1346.660 635.600 ;
      RECT 1348.620 1.400 1348.900 635.600 ;
      RECT 1350.860 1.400 1351.140 635.600 ;
      RECT 1353.100 1.400 1353.380 635.600 ;
      RECT 1355.340 1.400 1355.620 635.600 ;
      RECT 1357.580 1.400 1357.860 635.600 ;
      RECT 1359.820 1.400 1360.100 635.600 ;
      RECT 1362.060 1.400 1362.340 635.600 ;
      RECT 1364.300 1.400 1364.580 635.600 ;
      RECT 1366.540 1.400 1366.820 635.600 ;
      RECT 1368.780 1.400 1369.060 635.600 ;
      RECT 1371.020 1.400 1371.300 635.600 ;
      RECT 1373.260 1.400 1373.540 635.600 ;
      RECT 1375.500 1.400 1375.780 635.600 ;
      RECT 1377.740 1.400 1378.020 635.600 ;
      RECT 1379.980 1.400 1380.260 635.600 ;
      RECT 1382.220 1.400 1382.500 635.600 ;
      RECT 1384.460 1.400 1384.740 635.600 ;
      RECT 1386.700 1.400 1386.980 635.600 ;
      RECT 1388.940 1.400 1389.220 635.600 ;
      RECT 1391.180 1.400 1391.460 635.600 ;
      RECT 1393.420 1.400 1393.700 635.600 ;
      RECT 1395.660 1.400 1395.940 635.600 ;
      RECT 1397.900 1.400 1398.180 635.600 ;
      RECT 1400.140 1.400 1400.420 635.600 ;
      RECT 1402.380 1.400 1402.660 635.600 ;
      RECT 1404.620 1.400 1404.900 635.600 ;
      RECT 1406.860 1.400 1407.140 635.600 ;
      RECT 1409.100 1.400 1409.380 635.600 ;
      RECT 1411.340 1.400 1411.620 635.600 ;
      RECT 1413.580 1.400 1413.860 635.600 ;
      RECT 1415.820 1.400 1416.100 635.600 ;
      RECT 1418.060 1.400 1418.340 635.600 ;
      RECT 1420.300 1.400 1420.580 635.600 ;
      RECT 1422.540 1.400 1422.820 635.600 ;
      RECT 1424.780 1.400 1425.060 635.600 ;
      RECT 1427.020 1.400 1427.300 635.600 ;
      RECT 1429.260 1.400 1429.540 635.600 ;
      RECT 1431.500 1.400 1431.780 635.600 ;
      RECT 1433.740 1.400 1434.020 635.600 ;
      RECT 1435.980 1.400 1436.260 635.600 ;
      RECT 1438.220 1.400 1438.500 635.600 ;
      RECT 1440.460 1.400 1440.740 635.600 ;
      RECT 1442.700 1.400 1442.980 635.600 ;
      RECT 1444.940 1.400 1445.220 635.600 ;
      RECT 1447.180 1.400 1447.460 635.600 ;
      RECT 1449.420 1.400 1449.700 635.600 ;
      RECT 1451.660 1.400 1451.940 635.600 ;
      RECT 1453.900 1.400 1454.180 635.600 ;
      RECT 1456.140 1.400 1456.420 635.600 ;
      RECT 1458.380 1.400 1458.660 635.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 1461.480 637.000 ;
    LAYER metal2 ;
    RECT 0 0 1461.480 637.000 ;
    LAYER metal3 ;
    RECT 0.070 0 1461.480 637.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 4.305 ;
    RECT 0 4.375 0.070 7.245 ;
    RECT 0 7.315 0.070 10.185 ;
    RECT 0 10.255 0.070 13.125 ;
    RECT 0 13.195 0.070 16.065 ;
    RECT 0 16.135 0.070 19.005 ;
    RECT 0 19.075 0.070 21.945 ;
    RECT 0 22.015 0.070 24.885 ;
    RECT 0 24.955 0.070 27.825 ;
    RECT 0 27.895 0.070 30.765 ;
    RECT 0 30.835 0.070 33.705 ;
    RECT 0 33.775 0.070 36.645 ;
    RECT 0 36.715 0.070 39.585 ;
    RECT 0 39.655 0.070 42.525 ;
    RECT 0 42.595 0.070 45.465 ;
    RECT 0 45.535 0.070 48.405 ;
    RECT 0 48.475 0.070 51.345 ;
    RECT 0 51.415 0.070 54.285 ;
    RECT 0 54.355 0.070 57.225 ;
    RECT 0 57.295 0.070 60.165 ;
    RECT 0 60.235 0.070 63.105 ;
    RECT 0 63.175 0.070 66.045 ;
    RECT 0 66.115 0.070 68.985 ;
    RECT 0 69.055 0.070 71.925 ;
    RECT 0 71.995 0.070 74.865 ;
    RECT 0 74.935 0.070 77.805 ;
    RECT 0 77.875 0.070 80.745 ;
    RECT 0 80.815 0.070 83.685 ;
    RECT 0 83.755 0.070 86.625 ;
    RECT 0 86.695 0.070 89.565 ;
    RECT 0 89.635 0.070 92.505 ;
    RECT 0 92.575 0.070 95.445 ;
    RECT 0 95.515 0.070 98.385 ;
    RECT 0 98.455 0.070 101.325 ;
    RECT 0 101.395 0.070 104.265 ;
    RECT 0 104.335 0.070 107.205 ;
    RECT 0 107.275 0.070 110.145 ;
    RECT 0 110.215 0.070 113.085 ;
    RECT 0 113.155 0.070 116.025 ;
    RECT 0 116.095 0.070 118.965 ;
    RECT 0 119.035 0.070 121.905 ;
    RECT 0 121.975 0.070 124.845 ;
    RECT 0 124.915 0.070 127.785 ;
    RECT 0 127.855 0.070 130.725 ;
    RECT 0 130.795 0.070 133.665 ;
    RECT 0 133.735 0.070 136.605 ;
    RECT 0 136.675 0.070 139.545 ;
    RECT 0 139.615 0.070 142.485 ;
    RECT 0 142.555 0.070 145.425 ;
    RECT 0 145.495 0.070 148.365 ;
    RECT 0 148.435 0.070 151.305 ;
    RECT 0 151.375 0.070 154.245 ;
    RECT 0 154.315 0.070 157.185 ;
    RECT 0 157.255 0.070 160.125 ;
    RECT 0 160.195 0.070 163.065 ;
    RECT 0 163.135 0.070 166.005 ;
    RECT 0 166.075 0.070 168.945 ;
    RECT 0 169.015 0.070 171.885 ;
    RECT 0 171.955 0.070 174.825 ;
    RECT 0 174.895 0.070 177.765 ;
    RECT 0 177.835 0.070 180.705 ;
    RECT 0 180.775 0.070 183.645 ;
    RECT 0 183.715 0.070 186.585 ;
    RECT 0 186.655 0.070 191.485 ;
    RECT 0 191.555 0.070 194.425 ;
    RECT 0 194.495 0.070 197.365 ;
    RECT 0 197.435 0.070 200.305 ;
    RECT 0 200.375 0.070 203.245 ;
    RECT 0 203.315 0.070 206.185 ;
    RECT 0 206.255 0.070 209.125 ;
    RECT 0 209.195 0.070 212.065 ;
    RECT 0 212.135 0.070 215.005 ;
    RECT 0 215.075 0.070 217.945 ;
    RECT 0 218.015 0.070 220.885 ;
    RECT 0 220.955 0.070 223.825 ;
    RECT 0 223.895 0.070 226.765 ;
    RECT 0 226.835 0.070 229.705 ;
    RECT 0 229.775 0.070 232.645 ;
    RECT 0 232.715 0.070 235.585 ;
    RECT 0 235.655 0.070 238.525 ;
    RECT 0 238.595 0.070 241.465 ;
    RECT 0 241.535 0.070 244.405 ;
    RECT 0 244.475 0.070 247.345 ;
    RECT 0 247.415 0.070 250.285 ;
    RECT 0 250.355 0.070 253.225 ;
    RECT 0 253.295 0.070 256.165 ;
    RECT 0 256.235 0.070 259.105 ;
    RECT 0 259.175 0.070 262.045 ;
    RECT 0 262.115 0.070 264.985 ;
    RECT 0 265.055 0.070 267.925 ;
    RECT 0 267.995 0.070 270.865 ;
    RECT 0 270.935 0.070 273.805 ;
    RECT 0 273.875 0.070 276.745 ;
    RECT 0 276.815 0.070 279.685 ;
    RECT 0 279.755 0.070 282.625 ;
    RECT 0 282.695 0.070 285.565 ;
    RECT 0 285.635 0.070 288.505 ;
    RECT 0 288.575 0.070 291.445 ;
    RECT 0 291.515 0.070 294.385 ;
    RECT 0 294.455 0.070 297.325 ;
    RECT 0 297.395 0.070 300.265 ;
    RECT 0 300.335 0.070 303.205 ;
    RECT 0 303.275 0.070 306.145 ;
    RECT 0 306.215 0.070 309.085 ;
    RECT 0 309.155 0.070 312.025 ;
    RECT 0 312.095 0.070 314.965 ;
    RECT 0 315.035 0.070 317.905 ;
    RECT 0 317.975 0.070 320.845 ;
    RECT 0 320.915 0.070 323.785 ;
    RECT 0 323.855 0.070 326.725 ;
    RECT 0 326.795 0.070 329.665 ;
    RECT 0 329.735 0.070 332.605 ;
    RECT 0 332.675 0.070 335.545 ;
    RECT 0 335.615 0.070 338.485 ;
    RECT 0 338.555 0.070 341.425 ;
    RECT 0 341.495 0.070 344.365 ;
    RECT 0 344.435 0.070 347.305 ;
    RECT 0 347.375 0.070 350.245 ;
    RECT 0 350.315 0.070 353.185 ;
    RECT 0 353.255 0.070 356.125 ;
    RECT 0 356.195 0.070 359.065 ;
    RECT 0 359.135 0.070 362.005 ;
    RECT 0 362.075 0.070 364.945 ;
    RECT 0 365.015 0.070 367.885 ;
    RECT 0 367.955 0.070 370.825 ;
    RECT 0 370.895 0.070 373.765 ;
    RECT 0 373.835 0.070 376.705 ;
    RECT 0 376.775 0.070 381.605 ;
    RECT 0 381.675 0.070 384.545 ;
    RECT 0 384.615 0.070 387.485 ;
    RECT 0 387.555 0.070 390.425 ;
    RECT 0 390.495 0.070 393.365 ;
    RECT 0 393.435 0.070 396.305 ;
    RECT 0 396.375 0.070 399.245 ;
    RECT 0 399.315 0.070 402.185 ;
    RECT 0 402.255 0.070 405.125 ;
    RECT 0 405.195 0.070 408.065 ;
    RECT 0 408.135 0.070 411.005 ;
    RECT 0 411.075 0.070 413.945 ;
    RECT 0 414.015 0.070 416.885 ;
    RECT 0 416.955 0.070 419.825 ;
    RECT 0 419.895 0.070 422.765 ;
    RECT 0 422.835 0.070 425.705 ;
    RECT 0 425.775 0.070 428.645 ;
    RECT 0 428.715 0.070 431.585 ;
    RECT 0 431.655 0.070 434.525 ;
    RECT 0 434.595 0.070 437.465 ;
    RECT 0 437.535 0.070 440.405 ;
    RECT 0 440.475 0.070 443.345 ;
    RECT 0 443.415 0.070 446.285 ;
    RECT 0 446.355 0.070 449.225 ;
    RECT 0 449.295 0.070 452.165 ;
    RECT 0 452.235 0.070 455.105 ;
    RECT 0 455.175 0.070 458.045 ;
    RECT 0 458.115 0.070 460.985 ;
    RECT 0 461.055 0.070 463.925 ;
    RECT 0 463.995 0.070 466.865 ;
    RECT 0 466.935 0.070 469.805 ;
    RECT 0 469.875 0.070 472.745 ;
    RECT 0 472.815 0.070 475.685 ;
    RECT 0 475.755 0.070 478.625 ;
    RECT 0 478.695 0.070 481.565 ;
    RECT 0 481.635 0.070 484.505 ;
    RECT 0 484.575 0.070 487.445 ;
    RECT 0 487.515 0.070 490.385 ;
    RECT 0 490.455 0.070 493.325 ;
    RECT 0 493.395 0.070 496.265 ;
    RECT 0 496.335 0.070 499.205 ;
    RECT 0 499.275 0.070 502.145 ;
    RECT 0 502.215 0.070 505.085 ;
    RECT 0 505.155 0.070 508.025 ;
    RECT 0 508.095 0.070 510.965 ;
    RECT 0 511.035 0.070 513.905 ;
    RECT 0 513.975 0.070 516.845 ;
    RECT 0 516.915 0.070 519.785 ;
    RECT 0 519.855 0.070 522.725 ;
    RECT 0 522.795 0.070 525.665 ;
    RECT 0 525.735 0.070 528.605 ;
    RECT 0 528.675 0.070 531.545 ;
    RECT 0 531.615 0.070 534.485 ;
    RECT 0 534.555 0.070 537.425 ;
    RECT 0 537.495 0.070 540.365 ;
    RECT 0 540.435 0.070 543.305 ;
    RECT 0 543.375 0.070 546.245 ;
    RECT 0 546.315 0.070 549.185 ;
    RECT 0 549.255 0.070 552.125 ;
    RECT 0 552.195 0.070 555.065 ;
    RECT 0 555.135 0.070 558.005 ;
    RECT 0 558.075 0.070 560.945 ;
    RECT 0 561.015 0.070 563.885 ;
    RECT 0 563.955 0.070 566.825 ;
    RECT 0 566.895 0.070 571.725 ;
    RECT 0 571.795 0.070 574.665 ;
    RECT 0 574.735 0.070 577.605 ;
    RECT 0 577.675 0.070 580.545 ;
    RECT 0 580.615 0.070 583.485 ;
    RECT 0 583.555 0.070 586.425 ;
    RECT 0 586.495 0.070 589.365 ;
    RECT 0 589.435 0.070 592.305 ;
    RECT 0 592.375 0.070 595.245 ;
    RECT 0 595.315 0.070 598.185 ;
    RECT 0 598.255 0.070 601.125 ;
    RECT 0 601.195 0.070 604.065 ;
    RECT 0 604.135 0.070 607.005 ;
    RECT 0 607.075 0.070 609.945 ;
    RECT 0 610.015 0.070 614.845 ;
    RECT 0 614.915 0.070 617.785 ;
    RECT 0 617.855 0.070 620.725 ;
    RECT 0 620.795 0.070 637.000 ;
    LAYER metal4 ;
    RECT 0 0 1461.480 1.400 ;
    RECT 0 635.600 1461.480 637.000 ;
    RECT 0.000 1.400 1.260 635.600 ;
    RECT 1.540 1.400 2.380 635.600 ;
    RECT 2.660 1.400 3.500 635.600 ;
    RECT 3.780 1.400 4.620 635.600 ;
    RECT 4.900 1.400 5.740 635.600 ;
    RECT 6.020 1.400 6.860 635.600 ;
    RECT 7.140 1.400 7.980 635.600 ;
    RECT 8.260 1.400 9.100 635.600 ;
    RECT 9.380 1.400 10.220 635.600 ;
    RECT 10.500 1.400 11.340 635.600 ;
    RECT 11.620 1.400 12.460 635.600 ;
    RECT 12.740 1.400 13.580 635.600 ;
    RECT 13.860 1.400 14.700 635.600 ;
    RECT 14.980 1.400 15.820 635.600 ;
    RECT 16.100 1.400 16.940 635.600 ;
    RECT 17.220 1.400 18.060 635.600 ;
    RECT 18.340 1.400 19.180 635.600 ;
    RECT 19.460 1.400 20.300 635.600 ;
    RECT 20.580 1.400 21.420 635.600 ;
    RECT 21.700 1.400 22.540 635.600 ;
    RECT 22.820 1.400 23.660 635.600 ;
    RECT 23.940 1.400 24.780 635.600 ;
    RECT 25.060 1.400 25.900 635.600 ;
    RECT 26.180 1.400 27.020 635.600 ;
    RECT 27.300 1.400 28.140 635.600 ;
    RECT 28.420 1.400 29.260 635.600 ;
    RECT 29.540 1.400 30.380 635.600 ;
    RECT 30.660 1.400 31.500 635.600 ;
    RECT 31.780 1.400 32.620 635.600 ;
    RECT 32.900 1.400 33.740 635.600 ;
    RECT 34.020 1.400 34.860 635.600 ;
    RECT 35.140 1.400 35.980 635.600 ;
    RECT 36.260 1.400 37.100 635.600 ;
    RECT 37.380 1.400 38.220 635.600 ;
    RECT 38.500 1.400 39.340 635.600 ;
    RECT 39.620 1.400 40.460 635.600 ;
    RECT 40.740 1.400 41.580 635.600 ;
    RECT 41.860 1.400 42.700 635.600 ;
    RECT 42.980 1.400 43.820 635.600 ;
    RECT 44.100 1.400 44.940 635.600 ;
    RECT 45.220 1.400 46.060 635.600 ;
    RECT 46.340 1.400 47.180 635.600 ;
    RECT 47.460 1.400 48.300 635.600 ;
    RECT 48.580 1.400 49.420 635.600 ;
    RECT 49.700 1.400 50.540 635.600 ;
    RECT 50.820 1.400 51.660 635.600 ;
    RECT 51.940 1.400 52.780 635.600 ;
    RECT 53.060 1.400 53.900 635.600 ;
    RECT 54.180 1.400 55.020 635.600 ;
    RECT 55.300 1.400 56.140 635.600 ;
    RECT 56.420 1.400 57.260 635.600 ;
    RECT 57.540 1.400 58.380 635.600 ;
    RECT 58.660 1.400 59.500 635.600 ;
    RECT 59.780 1.400 60.620 635.600 ;
    RECT 60.900 1.400 61.740 635.600 ;
    RECT 62.020 1.400 62.860 635.600 ;
    RECT 63.140 1.400 63.980 635.600 ;
    RECT 64.260 1.400 65.100 635.600 ;
    RECT 65.380 1.400 66.220 635.600 ;
    RECT 66.500 1.400 67.340 635.600 ;
    RECT 67.620 1.400 68.460 635.600 ;
    RECT 68.740 1.400 69.580 635.600 ;
    RECT 69.860 1.400 70.700 635.600 ;
    RECT 70.980 1.400 71.820 635.600 ;
    RECT 72.100 1.400 72.940 635.600 ;
    RECT 73.220 1.400 74.060 635.600 ;
    RECT 74.340 1.400 75.180 635.600 ;
    RECT 75.460 1.400 76.300 635.600 ;
    RECT 76.580 1.400 77.420 635.600 ;
    RECT 77.700 1.400 78.540 635.600 ;
    RECT 78.820 1.400 79.660 635.600 ;
    RECT 79.940 1.400 80.780 635.600 ;
    RECT 81.060 1.400 81.900 635.600 ;
    RECT 82.180 1.400 83.020 635.600 ;
    RECT 83.300 1.400 84.140 635.600 ;
    RECT 84.420 1.400 85.260 635.600 ;
    RECT 85.540 1.400 86.380 635.600 ;
    RECT 86.660 1.400 87.500 635.600 ;
    RECT 87.780 1.400 88.620 635.600 ;
    RECT 88.900 1.400 89.740 635.600 ;
    RECT 90.020 1.400 90.860 635.600 ;
    RECT 91.140 1.400 91.980 635.600 ;
    RECT 92.260 1.400 93.100 635.600 ;
    RECT 93.380 1.400 94.220 635.600 ;
    RECT 94.500 1.400 95.340 635.600 ;
    RECT 95.620 1.400 96.460 635.600 ;
    RECT 96.740 1.400 97.580 635.600 ;
    RECT 97.860 1.400 98.700 635.600 ;
    RECT 98.980 1.400 99.820 635.600 ;
    RECT 100.100 1.400 100.940 635.600 ;
    RECT 101.220 1.400 102.060 635.600 ;
    RECT 102.340 1.400 103.180 635.600 ;
    RECT 103.460 1.400 104.300 635.600 ;
    RECT 104.580 1.400 105.420 635.600 ;
    RECT 105.700 1.400 106.540 635.600 ;
    RECT 106.820 1.400 107.660 635.600 ;
    RECT 107.940 1.400 108.780 635.600 ;
    RECT 109.060 1.400 109.900 635.600 ;
    RECT 110.180 1.400 111.020 635.600 ;
    RECT 111.300 1.400 112.140 635.600 ;
    RECT 112.420 1.400 113.260 635.600 ;
    RECT 113.540 1.400 114.380 635.600 ;
    RECT 114.660 1.400 115.500 635.600 ;
    RECT 115.780 1.400 116.620 635.600 ;
    RECT 116.900 1.400 117.740 635.600 ;
    RECT 118.020 1.400 118.860 635.600 ;
    RECT 119.140 1.400 119.980 635.600 ;
    RECT 120.260 1.400 121.100 635.600 ;
    RECT 121.380 1.400 122.220 635.600 ;
    RECT 122.500 1.400 123.340 635.600 ;
    RECT 123.620 1.400 124.460 635.600 ;
    RECT 124.740 1.400 125.580 635.600 ;
    RECT 125.860 1.400 126.700 635.600 ;
    RECT 126.980 1.400 127.820 635.600 ;
    RECT 128.100 1.400 128.940 635.600 ;
    RECT 129.220 1.400 130.060 635.600 ;
    RECT 130.340 1.400 131.180 635.600 ;
    RECT 131.460 1.400 132.300 635.600 ;
    RECT 132.580 1.400 133.420 635.600 ;
    RECT 133.700 1.400 134.540 635.600 ;
    RECT 134.820 1.400 135.660 635.600 ;
    RECT 135.940 1.400 136.780 635.600 ;
    RECT 137.060 1.400 137.900 635.600 ;
    RECT 138.180 1.400 139.020 635.600 ;
    RECT 139.300 1.400 140.140 635.600 ;
    RECT 140.420 1.400 141.260 635.600 ;
    RECT 141.540 1.400 142.380 635.600 ;
    RECT 142.660 1.400 143.500 635.600 ;
    RECT 143.780 1.400 144.620 635.600 ;
    RECT 144.900 1.400 145.740 635.600 ;
    RECT 146.020 1.400 146.860 635.600 ;
    RECT 147.140 1.400 147.980 635.600 ;
    RECT 148.260 1.400 149.100 635.600 ;
    RECT 149.380 1.400 150.220 635.600 ;
    RECT 150.500 1.400 151.340 635.600 ;
    RECT 151.620 1.400 152.460 635.600 ;
    RECT 152.740 1.400 153.580 635.600 ;
    RECT 153.860 1.400 154.700 635.600 ;
    RECT 154.980 1.400 155.820 635.600 ;
    RECT 156.100 1.400 156.940 635.600 ;
    RECT 157.220 1.400 158.060 635.600 ;
    RECT 158.340 1.400 159.180 635.600 ;
    RECT 159.460 1.400 160.300 635.600 ;
    RECT 160.580 1.400 161.420 635.600 ;
    RECT 161.700 1.400 162.540 635.600 ;
    RECT 162.820 1.400 163.660 635.600 ;
    RECT 163.940 1.400 164.780 635.600 ;
    RECT 165.060 1.400 165.900 635.600 ;
    RECT 166.180 1.400 167.020 635.600 ;
    RECT 167.300 1.400 168.140 635.600 ;
    RECT 168.420 1.400 169.260 635.600 ;
    RECT 169.540 1.400 170.380 635.600 ;
    RECT 170.660 1.400 171.500 635.600 ;
    RECT 171.780 1.400 172.620 635.600 ;
    RECT 172.900 1.400 173.740 635.600 ;
    RECT 174.020 1.400 174.860 635.600 ;
    RECT 175.140 1.400 175.980 635.600 ;
    RECT 176.260 1.400 177.100 635.600 ;
    RECT 177.380 1.400 178.220 635.600 ;
    RECT 178.500 1.400 179.340 635.600 ;
    RECT 179.620 1.400 180.460 635.600 ;
    RECT 180.740 1.400 181.580 635.600 ;
    RECT 181.860 1.400 182.700 635.600 ;
    RECT 182.980 1.400 183.820 635.600 ;
    RECT 184.100 1.400 184.940 635.600 ;
    RECT 185.220 1.400 186.060 635.600 ;
    RECT 186.340 1.400 187.180 635.600 ;
    RECT 187.460 1.400 188.300 635.600 ;
    RECT 188.580 1.400 189.420 635.600 ;
    RECT 189.700 1.400 190.540 635.600 ;
    RECT 190.820 1.400 191.660 635.600 ;
    RECT 191.940 1.400 192.780 635.600 ;
    RECT 193.060 1.400 193.900 635.600 ;
    RECT 194.180 1.400 195.020 635.600 ;
    RECT 195.300 1.400 196.140 635.600 ;
    RECT 196.420 1.400 197.260 635.600 ;
    RECT 197.540 1.400 198.380 635.600 ;
    RECT 198.660 1.400 199.500 635.600 ;
    RECT 199.780 1.400 200.620 635.600 ;
    RECT 200.900 1.400 201.740 635.600 ;
    RECT 202.020 1.400 202.860 635.600 ;
    RECT 203.140 1.400 203.980 635.600 ;
    RECT 204.260 1.400 205.100 635.600 ;
    RECT 205.380 1.400 206.220 635.600 ;
    RECT 206.500 1.400 207.340 635.600 ;
    RECT 207.620 1.400 208.460 635.600 ;
    RECT 208.740 1.400 209.580 635.600 ;
    RECT 209.860 1.400 210.700 635.600 ;
    RECT 210.980 1.400 211.820 635.600 ;
    RECT 212.100 1.400 212.940 635.600 ;
    RECT 213.220 1.400 214.060 635.600 ;
    RECT 214.340 1.400 215.180 635.600 ;
    RECT 215.460 1.400 216.300 635.600 ;
    RECT 216.580 1.400 217.420 635.600 ;
    RECT 217.700 1.400 218.540 635.600 ;
    RECT 218.820 1.400 219.660 635.600 ;
    RECT 219.940 1.400 220.780 635.600 ;
    RECT 221.060 1.400 221.900 635.600 ;
    RECT 222.180 1.400 223.020 635.600 ;
    RECT 223.300 1.400 224.140 635.600 ;
    RECT 224.420 1.400 225.260 635.600 ;
    RECT 225.540 1.400 226.380 635.600 ;
    RECT 226.660 1.400 227.500 635.600 ;
    RECT 227.780 1.400 228.620 635.600 ;
    RECT 228.900 1.400 229.740 635.600 ;
    RECT 230.020 1.400 230.860 635.600 ;
    RECT 231.140 1.400 231.980 635.600 ;
    RECT 232.260 1.400 233.100 635.600 ;
    RECT 233.380 1.400 234.220 635.600 ;
    RECT 234.500 1.400 235.340 635.600 ;
    RECT 235.620 1.400 236.460 635.600 ;
    RECT 236.740 1.400 237.580 635.600 ;
    RECT 237.860 1.400 238.700 635.600 ;
    RECT 238.980 1.400 239.820 635.600 ;
    RECT 240.100 1.400 240.940 635.600 ;
    RECT 241.220 1.400 242.060 635.600 ;
    RECT 242.340 1.400 243.180 635.600 ;
    RECT 243.460 1.400 244.300 635.600 ;
    RECT 244.580 1.400 245.420 635.600 ;
    RECT 245.700 1.400 246.540 635.600 ;
    RECT 246.820 1.400 247.660 635.600 ;
    RECT 247.940 1.400 248.780 635.600 ;
    RECT 249.060 1.400 249.900 635.600 ;
    RECT 250.180 1.400 251.020 635.600 ;
    RECT 251.300 1.400 252.140 635.600 ;
    RECT 252.420 1.400 253.260 635.600 ;
    RECT 253.540 1.400 254.380 635.600 ;
    RECT 254.660 1.400 255.500 635.600 ;
    RECT 255.780 1.400 256.620 635.600 ;
    RECT 256.900 1.400 257.740 635.600 ;
    RECT 258.020 1.400 258.860 635.600 ;
    RECT 259.140 1.400 259.980 635.600 ;
    RECT 260.260 1.400 261.100 635.600 ;
    RECT 261.380 1.400 262.220 635.600 ;
    RECT 262.500 1.400 263.340 635.600 ;
    RECT 263.620 1.400 264.460 635.600 ;
    RECT 264.740 1.400 265.580 635.600 ;
    RECT 265.860 1.400 266.700 635.600 ;
    RECT 266.980 1.400 267.820 635.600 ;
    RECT 268.100 1.400 268.940 635.600 ;
    RECT 269.220 1.400 270.060 635.600 ;
    RECT 270.340 1.400 271.180 635.600 ;
    RECT 271.460 1.400 272.300 635.600 ;
    RECT 272.580 1.400 273.420 635.600 ;
    RECT 273.700 1.400 274.540 635.600 ;
    RECT 274.820 1.400 275.660 635.600 ;
    RECT 275.940 1.400 276.780 635.600 ;
    RECT 277.060 1.400 277.900 635.600 ;
    RECT 278.180 1.400 279.020 635.600 ;
    RECT 279.300 1.400 280.140 635.600 ;
    RECT 280.420 1.400 281.260 635.600 ;
    RECT 281.540 1.400 282.380 635.600 ;
    RECT 282.660 1.400 283.500 635.600 ;
    RECT 283.780 1.400 284.620 635.600 ;
    RECT 284.900 1.400 285.740 635.600 ;
    RECT 286.020 1.400 286.860 635.600 ;
    RECT 287.140 1.400 287.980 635.600 ;
    RECT 288.260 1.400 289.100 635.600 ;
    RECT 289.380 1.400 290.220 635.600 ;
    RECT 290.500 1.400 291.340 635.600 ;
    RECT 291.620 1.400 292.460 635.600 ;
    RECT 292.740 1.400 293.580 635.600 ;
    RECT 293.860 1.400 294.700 635.600 ;
    RECT 294.980 1.400 295.820 635.600 ;
    RECT 296.100 1.400 296.940 635.600 ;
    RECT 297.220 1.400 298.060 635.600 ;
    RECT 298.340 1.400 299.180 635.600 ;
    RECT 299.460 1.400 300.300 635.600 ;
    RECT 300.580 1.400 301.420 635.600 ;
    RECT 301.700 1.400 302.540 635.600 ;
    RECT 302.820 1.400 303.660 635.600 ;
    RECT 303.940 1.400 304.780 635.600 ;
    RECT 305.060 1.400 305.900 635.600 ;
    RECT 306.180 1.400 307.020 635.600 ;
    RECT 307.300 1.400 308.140 635.600 ;
    RECT 308.420 1.400 309.260 635.600 ;
    RECT 309.540 1.400 310.380 635.600 ;
    RECT 310.660 1.400 311.500 635.600 ;
    RECT 311.780 1.400 312.620 635.600 ;
    RECT 312.900 1.400 313.740 635.600 ;
    RECT 314.020 1.400 314.860 635.600 ;
    RECT 315.140 1.400 315.980 635.600 ;
    RECT 316.260 1.400 317.100 635.600 ;
    RECT 317.380 1.400 318.220 635.600 ;
    RECT 318.500 1.400 319.340 635.600 ;
    RECT 319.620 1.400 320.460 635.600 ;
    RECT 320.740 1.400 321.580 635.600 ;
    RECT 321.860 1.400 322.700 635.600 ;
    RECT 322.980 1.400 323.820 635.600 ;
    RECT 324.100 1.400 324.940 635.600 ;
    RECT 325.220 1.400 326.060 635.600 ;
    RECT 326.340 1.400 327.180 635.600 ;
    RECT 327.460 1.400 328.300 635.600 ;
    RECT 328.580 1.400 329.420 635.600 ;
    RECT 329.700 1.400 330.540 635.600 ;
    RECT 330.820 1.400 331.660 635.600 ;
    RECT 331.940 1.400 332.780 635.600 ;
    RECT 333.060 1.400 333.900 635.600 ;
    RECT 334.180 1.400 335.020 635.600 ;
    RECT 335.300 1.400 336.140 635.600 ;
    RECT 336.420 1.400 337.260 635.600 ;
    RECT 337.540 1.400 338.380 635.600 ;
    RECT 338.660 1.400 339.500 635.600 ;
    RECT 339.780 1.400 340.620 635.600 ;
    RECT 340.900 1.400 341.740 635.600 ;
    RECT 342.020 1.400 342.860 635.600 ;
    RECT 343.140 1.400 343.980 635.600 ;
    RECT 344.260 1.400 345.100 635.600 ;
    RECT 345.380 1.400 346.220 635.600 ;
    RECT 346.500 1.400 347.340 635.600 ;
    RECT 347.620 1.400 348.460 635.600 ;
    RECT 348.740 1.400 349.580 635.600 ;
    RECT 349.860 1.400 350.700 635.600 ;
    RECT 350.980 1.400 351.820 635.600 ;
    RECT 352.100 1.400 352.940 635.600 ;
    RECT 353.220 1.400 354.060 635.600 ;
    RECT 354.340 1.400 355.180 635.600 ;
    RECT 355.460 1.400 356.300 635.600 ;
    RECT 356.580 1.400 357.420 635.600 ;
    RECT 357.700 1.400 358.540 635.600 ;
    RECT 358.820 1.400 359.660 635.600 ;
    RECT 359.940 1.400 360.780 635.600 ;
    RECT 361.060 1.400 361.900 635.600 ;
    RECT 362.180 1.400 363.020 635.600 ;
    RECT 363.300 1.400 364.140 635.600 ;
    RECT 364.420 1.400 365.260 635.600 ;
    RECT 365.540 1.400 366.380 635.600 ;
    RECT 366.660 1.400 367.500 635.600 ;
    RECT 367.780 1.400 368.620 635.600 ;
    RECT 368.900 1.400 369.740 635.600 ;
    RECT 370.020 1.400 370.860 635.600 ;
    RECT 371.140 1.400 371.980 635.600 ;
    RECT 372.260 1.400 373.100 635.600 ;
    RECT 373.380 1.400 374.220 635.600 ;
    RECT 374.500 1.400 375.340 635.600 ;
    RECT 375.620 1.400 376.460 635.600 ;
    RECT 376.740 1.400 377.580 635.600 ;
    RECT 377.860 1.400 378.700 635.600 ;
    RECT 378.980 1.400 379.820 635.600 ;
    RECT 380.100 1.400 380.940 635.600 ;
    RECT 381.220 1.400 382.060 635.600 ;
    RECT 382.340 1.400 383.180 635.600 ;
    RECT 383.460 1.400 384.300 635.600 ;
    RECT 384.580 1.400 385.420 635.600 ;
    RECT 385.700 1.400 386.540 635.600 ;
    RECT 386.820 1.400 387.660 635.600 ;
    RECT 387.940 1.400 388.780 635.600 ;
    RECT 389.060 1.400 389.900 635.600 ;
    RECT 390.180 1.400 391.020 635.600 ;
    RECT 391.300 1.400 392.140 635.600 ;
    RECT 392.420 1.400 393.260 635.600 ;
    RECT 393.540 1.400 394.380 635.600 ;
    RECT 394.660 1.400 395.500 635.600 ;
    RECT 395.780 1.400 396.620 635.600 ;
    RECT 396.900 1.400 397.740 635.600 ;
    RECT 398.020 1.400 398.860 635.600 ;
    RECT 399.140 1.400 399.980 635.600 ;
    RECT 400.260 1.400 401.100 635.600 ;
    RECT 401.380 1.400 402.220 635.600 ;
    RECT 402.500 1.400 403.340 635.600 ;
    RECT 403.620 1.400 404.460 635.600 ;
    RECT 404.740 1.400 405.580 635.600 ;
    RECT 405.860 1.400 406.700 635.600 ;
    RECT 406.980 1.400 407.820 635.600 ;
    RECT 408.100 1.400 408.940 635.600 ;
    RECT 409.220 1.400 410.060 635.600 ;
    RECT 410.340 1.400 411.180 635.600 ;
    RECT 411.460 1.400 412.300 635.600 ;
    RECT 412.580 1.400 413.420 635.600 ;
    RECT 413.700 1.400 414.540 635.600 ;
    RECT 414.820 1.400 415.660 635.600 ;
    RECT 415.940 1.400 416.780 635.600 ;
    RECT 417.060 1.400 417.900 635.600 ;
    RECT 418.180 1.400 419.020 635.600 ;
    RECT 419.300 1.400 420.140 635.600 ;
    RECT 420.420 1.400 421.260 635.600 ;
    RECT 421.540 1.400 422.380 635.600 ;
    RECT 422.660 1.400 423.500 635.600 ;
    RECT 423.780 1.400 424.620 635.600 ;
    RECT 424.900 1.400 425.740 635.600 ;
    RECT 426.020 1.400 426.860 635.600 ;
    RECT 427.140 1.400 427.980 635.600 ;
    RECT 428.260 1.400 429.100 635.600 ;
    RECT 429.380 1.400 430.220 635.600 ;
    RECT 430.500 1.400 431.340 635.600 ;
    RECT 431.620 1.400 432.460 635.600 ;
    RECT 432.740 1.400 433.580 635.600 ;
    RECT 433.860 1.400 434.700 635.600 ;
    RECT 434.980 1.400 435.820 635.600 ;
    RECT 436.100 1.400 436.940 635.600 ;
    RECT 437.220 1.400 438.060 635.600 ;
    RECT 438.340 1.400 439.180 635.600 ;
    RECT 439.460 1.400 440.300 635.600 ;
    RECT 440.580 1.400 441.420 635.600 ;
    RECT 441.700 1.400 442.540 635.600 ;
    RECT 442.820 1.400 443.660 635.600 ;
    RECT 443.940 1.400 444.780 635.600 ;
    RECT 445.060 1.400 445.900 635.600 ;
    RECT 446.180 1.400 447.020 635.600 ;
    RECT 447.300 1.400 448.140 635.600 ;
    RECT 448.420 1.400 449.260 635.600 ;
    RECT 449.540 1.400 450.380 635.600 ;
    RECT 450.660 1.400 451.500 635.600 ;
    RECT 451.780 1.400 452.620 635.600 ;
    RECT 452.900 1.400 453.740 635.600 ;
    RECT 454.020 1.400 454.860 635.600 ;
    RECT 455.140 1.400 455.980 635.600 ;
    RECT 456.260 1.400 457.100 635.600 ;
    RECT 457.380 1.400 458.220 635.600 ;
    RECT 458.500 1.400 459.340 635.600 ;
    RECT 459.620 1.400 460.460 635.600 ;
    RECT 460.740 1.400 461.580 635.600 ;
    RECT 461.860 1.400 462.700 635.600 ;
    RECT 462.980 1.400 463.820 635.600 ;
    RECT 464.100 1.400 464.940 635.600 ;
    RECT 465.220 1.400 466.060 635.600 ;
    RECT 466.340 1.400 467.180 635.600 ;
    RECT 467.460 1.400 468.300 635.600 ;
    RECT 468.580 1.400 469.420 635.600 ;
    RECT 469.700 1.400 470.540 635.600 ;
    RECT 470.820 1.400 471.660 635.600 ;
    RECT 471.940 1.400 472.780 635.600 ;
    RECT 473.060 1.400 473.900 635.600 ;
    RECT 474.180 1.400 475.020 635.600 ;
    RECT 475.300 1.400 476.140 635.600 ;
    RECT 476.420 1.400 477.260 635.600 ;
    RECT 477.540 1.400 478.380 635.600 ;
    RECT 478.660 1.400 479.500 635.600 ;
    RECT 479.780 1.400 480.620 635.600 ;
    RECT 480.900 1.400 481.740 635.600 ;
    RECT 482.020 1.400 482.860 635.600 ;
    RECT 483.140 1.400 483.980 635.600 ;
    RECT 484.260 1.400 485.100 635.600 ;
    RECT 485.380 1.400 486.220 635.600 ;
    RECT 486.500 1.400 487.340 635.600 ;
    RECT 487.620 1.400 488.460 635.600 ;
    RECT 488.740 1.400 489.580 635.600 ;
    RECT 489.860 1.400 490.700 635.600 ;
    RECT 490.980 1.400 491.820 635.600 ;
    RECT 492.100 1.400 492.940 635.600 ;
    RECT 493.220 1.400 494.060 635.600 ;
    RECT 494.340 1.400 495.180 635.600 ;
    RECT 495.460 1.400 496.300 635.600 ;
    RECT 496.580 1.400 497.420 635.600 ;
    RECT 497.700 1.400 498.540 635.600 ;
    RECT 498.820 1.400 499.660 635.600 ;
    RECT 499.940 1.400 500.780 635.600 ;
    RECT 501.060 1.400 501.900 635.600 ;
    RECT 502.180 1.400 503.020 635.600 ;
    RECT 503.300 1.400 504.140 635.600 ;
    RECT 504.420 1.400 505.260 635.600 ;
    RECT 505.540 1.400 506.380 635.600 ;
    RECT 506.660 1.400 507.500 635.600 ;
    RECT 507.780 1.400 508.620 635.600 ;
    RECT 508.900 1.400 509.740 635.600 ;
    RECT 510.020 1.400 510.860 635.600 ;
    RECT 511.140 1.400 511.980 635.600 ;
    RECT 512.260 1.400 513.100 635.600 ;
    RECT 513.380 1.400 514.220 635.600 ;
    RECT 514.500 1.400 515.340 635.600 ;
    RECT 515.620 1.400 516.460 635.600 ;
    RECT 516.740 1.400 517.580 635.600 ;
    RECT 517.860 1.400 518.700 635.600 ;
    RECT 518.980 1.400 519.820 635.600 ;
    RECT 520.100 1.400 520.940 635.600 ;
    RECT 521.220 1.400 522.060 635.600 ;
    RECT 522.340 1.400 523.180 635.600 ;
    RECT 523.460 1.400 524.300 635.600 ;
    RECT 524.580 1.400 525.420 635.600 ;
    RECT 525.700 1.400 526.540 635.600 ;
    RECT 526.820 1.400 527.660 635.600 ;
    RECT 527.940 1.400 528.780 635.600 ;
    RECT 529.060 1.400 529.900 635.600 ;
    RECT 530.180 1.400 531.020 635.600 ;
    RECT 531.300 1.400 532.140 635.600 ;
    RECT 532.420 1.400 533.260 635.600 ;
    RECT 533.540 1.400 534.380 635.600 ;
    RECT 534.660 1.400 535.500 635.600 ;
    RECT 535.780 1.400 536.620 635.600 ;
    RECT 536.900 1.400 537.740 635.600 ;
    RECT 538.020 1.400 538.860 635.600 ;
    RECT 539.140 1.400 539.980 635.600 ;
    RECT 540.260 1.400 541.100 635.600 ;
    RECT 541.380 1.400 542.220 635.600 ;
    RECT 542.500 1.400 543.340 635.600 ;
    RECT 543.620 1.400 544.460 635.600 ;
    RECT 544.740 1.400 545.580 635.600 ;
    RECT 545.860 1.400 546.700 635.600 ;
    RECT 546.980 1.400 547.820 635.600 ;
    RECT 548.100 1.400 548.940 635.600 ;
    RECT 549.220 1.400 550.060 635.600 ;
    RECT 550.340 1.400 551.180 635.600 ;
    RECT 551.460 1.400 552.300 635.600 ;
    RECT 552.580 1.400 553.420 635.600 ;
    RECT 553.700 1.400 554.540 635.600 ;
    RECT 554.820 1.400 555.660 635.600 ;
    RECT 555.940 1.400 556.780 635.600 ;
    RECT 557.060 1.400 557.900 635.600 ;
    RECT 558.180 1.400 559.020 635.600 ;
    RECT 559.300 1.400 560.140 635.600 ;
    RECT 560.420 1.400 561.260 635.600 ;
    RECT 561.540 1.400 562.380 635.600 ;
    RECT 562.660 1.400 563.500 635.600 ;
    RECT 563.780 1.400 564.620 635.600 ;
    RECT 564.900 1.400 565.740 635.600 ;
    RECT 566.020 1.400 566.860 635.600 ;
    RECT 567.140 1.400 567.980 635.600 ;
    RECT 568.260 1.400 569.100 635.600 ;
    RECT 569.380 1.400 570.220 635.600 ;
    RECT 570.500 1.400 571.340 635.600 ;
    RECT 571.620 1.400 572.460 635.600 ;
    RECT 572.740 1.400 573.580 635.600 ;
    RECT 573.860 1.400 574.700 635.600 ;
    RECT 574.980 1.400 575.820 635.600 ;
    RECT 576.100 1.400 576.940 635.600 ;
    RECT 577.220 1.400 578.060 635.600 ;
    RECT 578.340 1.400 579.180 635.600 ;
    RECT 579.460 1.400 580.300 635.600 ;
    RECT 580.580 1.400 581.420 635.600 ;
    RECT 581.700 1.400 582.540 635.600 ;
    RECT 582.820 1.400 583.660 635.600 ;
    RECT 583.940 1.400 584.780 635.600 ;
    RECT 585.060 1.400 585.900 635.600 ;
    RECT 586.180 1.400 587.020 635.600 ;
    RECT 587.300 1.400 588.140 635.600 ;
    RECT 588.420 1.400 589.260 635.600 ;
    RECT 589.540 1.400 590.380 635.600 ;
    RECT 590.660 1.400 591.500 635.600 ;
    RECT 591.780 1.400 592.620 635.600 ;
    RECT 592.900 1.400 593.740 635.600 ;
    RECT 594.020 1.400 594.860 635.600 ;
    RECT 595.140 1.400 595.980 635.600 ;
    RECT 596.260 1.400 597.100 635.600 ;
    RECT 597.380 1.400 598.220 635.600 ;
    RECT 598.500 1.400 599.340 635.600 ;
    RECT 599.620 1.400 600.460 635.600 ;
    RECT 600.740 1.400 601.580 635.600 ;
    RECT 601.860 1.400 602.700 635.600 ;
    RECT 602.980 1.400 603.820 635.600 ;
    RECT 604.100 1.400 604.940 635.600 ;
    RECT 605.220 1.400 606.060 635.600 ;
    RECT 606.340 1.400 607.180 635.600 ;
    RECT 607.460 1.400 608.300 635.600 ;
    RECT 608.580 1.400 609.420 635.600 ;
    RECT 609.700 1.400 610.540 635.600 ;
    RECT 610.820 1.400 611.660 635.600 ;
    RECT 611.940 1.400 612.780 635.600 ;
    RECT 613.060 1.400 613.900 635.600 ;
    RECT 614.180 1.400 615.020 635.600 ;
    RECT 615.300 1.400 616.140 635.600 ;
    RECT 616.420 1.400 617.260 635.600 ;
    RECT 617.540 1.400 618.380 635.600 ;
    RECT 618.660 1.400 619.500 635.600 ;
    RECT 619.780 1.400 620.620 635.600 ;
    RECT 620.900 1.400 621.740 635.600 ;
    RECT 622.020 1.400 622.860 635.600 ;
    RECT 623.140 1.400 623.980 635.600 ;
    RECT 624.260 1.400 625.100 635.600 ;
    RECT 625.380 1.400 626.220 635.600 ;
    RECT 626.500 1.400 627.340 635.600 ;
    RECT 627.620 1.400 628.460 635.600 ;
    RECT 628.740 1.400 629.580 635.600 ;
    RECT 629.860 1.400 630.700 635.600 ;
    RECT 630.980 1.400 631.820 635.600 ;
    RECT 632.100 1.400 632.940 635.600 ;
    RECT 633.220 1.400 634.060 635.600 ;
    RECT 634.340 1.400 635.180 635.600 ;
    RECT 635.460 1.400 636.300 635.600 ;
    RECT 636.580 1.400 637.420 635.600 ;
    RECT 637.700 1.400 638.540 635.600 ;
    RECT 638.820 1.400 639.660 635.600 ;
    RECT 639.940 1.400 640.780 635.600 ;
    RECT 641.060 1.400 641.900 635.600 ;
    RECT 642.180 1.400 643.020 635.600 ;
    RECT 643.300 1.400 644.140 635.600 ;
    RECT 644.420 1.400 645.260 635.600 ;
    RECT 645.540 1.400 646.380 635.600 ;
    RECT 646.660 1.400 647.500 635.600 ;
    RECT 647.780 1.400 648.620 635.600 ;
    RECT 648.900 1.400 649.740 635.600 ;
    RECT 650.020 1.400 650.860 635.600 ;
    RECT 651.140 1.400 651.980 635.600 ;
    RECT 652.260 1.400 653.100 635.600 ;
    RECT 653.380 1.400 654.220 635.600 ;
    RECT 654.500 1.400 655.340 635.600 ;
    RECT 655.620 1.400 656.460 635.600 ;
    RECT 656.740 1.400 657.580 635.600 ;
    RECT 657.860 1.400 658.700 635.600 ;
    RECT 658.980 1.400 659.820 635.600 ;
    RECT 660.100 1.400 660.940 635.600 ;
    RECT 661.220 1.400 662.060 635.600 ;
    RECT 662.340 1.400 663.180 635.600 ;
    RECT 663.460 1.400 664.300 635.600 ;
    RECT 664.580 1.400 665.420 635.600 ;
    RECT 665.700 1.400 666.540 635.600 ;
    RECT 666.820 1.400 667.660 635.600 ;
    RECT 667.940 1.400 668.780 635.600 ;
    RECT 669.060 1.400 669.900 635.600 ;
    RECT 670.180 1.400 671.020 635.600 ;
    RECT 671.300 1.400 672.140 635.600 ;
    RECT 672.420 1.400 673.260 635.600 ;
    RECT 673.540 1.400 674.380 635.600 ;
    RECT 674.660 1.400 675.500 635.600 ;
    RECT 675.780 1.400 676.620 635.600 ;
    RECT 676.900 1.400 677.740 635.600 ;
    RECT 678.020 1.400 678.860 635.600 ;
    RECT 679.140 1.400 679.980 635.600 ;
    RECT 680.260 1.400 681.100 635.600 ;
    RECT 681.380 1.400 682.220 635.600 ;
    RECT 682.500 1.400 683.340 635.600 ;
    RECT 683.620 1.400 684.460 635.600 ;
    RECT 684.740 1.400 685.580 635.600 ;
    RECT 685.860 1.400 686.700 635.600 ;
    RECT 686.980 1.400 687.820 635.600 ;
    RECT 688.100 1.400 688.940 635.600 ;
    RECT 689.220 1.400 690.060 635.600 ;
    RECT 690.340 1.400 691.180 635.600 ;
    RECT 691.460 1.400 692.300 635.600 ;
    RECT 692.580 1.400 693.420 635.600 ;
    RECT 693.700 1.400 694.540 635.600 ;
    RECT 694.820 1.400 695.660 635.600 ;
    RECT 695.940 1.400 696.780 635.600 ;
    RECT 697.060 1.400 697.900 635.600 ;
    RECT 698.180 1.400 699.020 635.600 ;
    RECT 699.300 1.400 700.140 635.600 ;
    RECT 700.420 1.400 701.260 635.600 ;
    RECT 701.540 1.400 702.380 635.600 ;
    RECT 702.660 1.400 703.500 635.600 ;
    RECT 703.780 1.400 704.620 635.600 ;
    RECT 704.900 1.400 705.740 635.600 ;
    RECT 706.020 1.400 706.860 635.600 ;
    RECT 707.140 1.400 707.980 635.600 ;
    RECT 708.260 1.400 709.100 635.600 ;
    RECT 709.380 1.400 710.220 635.600 ;
    RECT 710.500 1.400 711.340 635.600 ;
    RECT 711.620 1.400 712.460 635.600 ;
    RECT 712.740 1.400 713.580 635.600 ;
    RECT 713.860 1.400 714.700 635.600 ;
    RECT 714.980 1.400 715.820 635.600 ;
    RECT 716.100 1.400 716.940 635.600 ;
    RECT 717.220 1.400 718.060 635.600 ;
    RECT 718.340 1.400 719.180 635.600 ;
    RECT 719.460 1.400 720.300 635.600 ;
    RECT 720.580 1.400 721.420 635.600 ;
    RECT 721.700 1.400 722.540 635.600 ;
    RECT 722.820 1.400 723.660 635.600 ;
    RECT 723.940 1.400 724.780 635.600 ;
    RECT 725.060 1.400 725.900 635.600 ;
    RECT 726.180 1.400 727.020 635.600 ;
    RECT 727.300 1.400 728.140 635.600 ;
    RECT 728.420 1.400 729.260 635.600 ;
    RECT 729.540 1.400 730.380 635.600 ;
    RECT 730.660 1.400 731.500 635.600 ;
    RECT 731.780 1.400 732.620 635.600 ;
    RECT 732.900 1.400 733.740 635.600 ;
    RECT 734.020 1.400 734.860 635.600 ;
    RECT 735.140 1.400 735.980 635.600 ;
    RECT 736.260 1.400 737.100 635.600 ;
    RECT 737.380 1.400 738.220 635.600 ;
    RECT 738.500 1.400 739.340 635.600 ;
    RECT 739.620 1.400 740.460 635.600 ;
    RECT 740.740 1.400 741.580 635.600 ;
    RECT 741.860 1.400 742.700 635.600 ;
    RECT 742.980 1.400 743.820 635.600 ;
    RECT 744.100 1.400 744.940 635.600 ;
    RECT 745.220 1.400 746.060 635.600 ;
    RECT 746.340 1.400 747.180 635.600 ;
    RECT 747.460 1.400 748.300 635.600 ;
    RECT 748.580 1.400 749.420 635.600 ;
    RECT 749.700 1.400 750.540 635.600 ;
    RECT 750.820 1.400 751.660 635.600 ;
    RECT 751.940 1.400 752.780 635.600 ;
    RECT 753.060 1.400 753.900 635.600 ;
    RECT 754.180 1.400 755.020 635.600 ;
    RECT 755.300 1.400 756.140 635.600 ;
    RECT 756.420 1.400 757.260 635.600 ;
    RECT 757.540 1.400 758.380 635.600 ;
    RECT 758.660 1.400 759.500 635.600 ;
    RECT 759.780 1.400 760.620 635.600 ;
    RECT 760.900 1.400 761.740 635.600 ;
    RECT 762.020 1.400 762.860 635.600 ;
    RECT 763.140 1.400 763.980 635.600 ;
    RECT 764.260 1.400 765.100 635.600 ;
    RECT 765.380 1.400 766.220 635.600 ;
    RECT 766.500 1.400 767.340 635.600 ;
    RECT 767.620 1.400 768.460 635.600 ;
    RECT 768.740 1.400 769.580 635.600 ;
    RECT 769.860 1.400 770.700 635.600 ;
    RECT 770.980 1.400 771.820 635.600 ;
    RECT 772.100 1.400 772.940 635.600 ;
    RECT 773.220 1.400 774.060 635.600 ;
    RECT 774.340 1.400 775.180 635.600 ;
    RECT 775.460 1.400 776.300 635.600 ;
    RECT 776.580 1.400 777.420 635.600 ;
    RECT 777.700 1.400 778.540 635.600 ;
    RECT 778.820 1.400 779.660 635.600 ;
    RECT 779.940 1.400 780.780 635.600 ;
    RECT 781.060 1.400 781.900 635.600 ;
    RECT 782.180 1.400 783.020 635.600 ;
    RECT 783.300 1.400 784.140 635.600 ;
    RECT 784.420 1.400 785.260 635.600 ;
    RECT 785.540 1.400 786.380 635.600 ;
    RECT 786.660 1.400 787.500 635.600 ;
    RECT 787.780 1.400 788.620 635.600 ;
    RECT 788.900 1.400 789.740 635.600 ;
    RECT 790.020 1.400 790.860 635.600 ;
    RECT 791.140 1.400 791.980 635.600 ;
    RECT 792.260 1.400 793.100 635.600 ;
    RECT 793.380 1.400 794.220 635.600 ;
    RECT 794.500 1.400 795.340 635.600 ;
    RECT 795.620 1.400 796.460 635.600 ;
    RECT 796.740 1.400 797.580 635.600 ;
    RECT 797.860 1.400 798.700 635.600 ;
    RECT 798.980 1.400 799.820 635.600 ;
    RECT 800.100 1.400 800.940 635.600 ;
    RECT 801.220 1.400 802.060 635.600 ;
    RECT 802.340 1.400 803.180 635.600 ;
    RECT 803.460 1.400 804.300 635.600 ;
    RECT 804.580 1.400 805.420 635.600 ;
    RECT 805.700 1.400 806.540 635.600 ;
    RECT 806.820 1.400 807.660 635.600 ;
    RECT 807.940 1.400 808.780 635.600 ;
    RECT 809.060 1.400 809.900 635.600 ;
    RECT 810.180 1.400 811.020 635.600 ;
    RECT 811.300 1.400 812.140 635.600 ;
    RECT 812.420 1.400 813.260 635.600 ;
    RECT 813.540 1.400 814.380 635.600 ;
    RECT 814.660 1.400 815.500 635.600 ;
    RECT 815.780 1.400 816.620 635.600 ;
    RECT 816.900 1.400 817.740 635.600 ;
    RECT 818.020 1.400 818.860 635.600 ;
    RECT 819.140 1.400 819.980 635.600 ;
    RECT 820.260 1.400 821.100 635.600 ;
    RECT 821.380 1.400 822.220 635.600 ;
    RECT 822.500 1.400 823.340 635.600 ;
    RECT 823.620 1.400 824.460 635.600 ;
    RECT 824.740 1.400 825.580 635.600 ;
    RECT 825.860 1.400 826.700 635.600 ;
    RECT 826.980 1.400 827.820 635.600 ;
    RECT 828.100 1.400 828.940 635.600 ;
    RECT 829.220 1.400 830.060 635.600 ;
    RECT 830.340 1.400 831.180 635.600 ;
    RECT 831.460 1.400 832.300 635.600 ;
    RECT 832.580 1.400 833.420 635.600 ;
    RECT 833.700 1.400 834.540 635.600 ;
    RECT 834.820 1.400 835.660 635.600 ;
    RECT 835.940 1.400 836.780 635.600 ;
    RECT 837.060 1.400 837.900 635.600 ;
    RECT 838.180 1.400 839.020 635.600 ;
    RECT 839.300 1.400 840.140 635.600 ;
    RECT 840.420 1.400 841.260 635.600 ;
    RECT 841.540 1.400 842.380 635.600 ;
    RECT 842.660 1.400 843.500 635.600 ;
    RECT 843.780 1.400 844.620 635.600 ;
    RECT 844.900 1.400 845.740 635.600 ;
    RECT 846.020 1.400 846.860 635.600 ;
    RECT 847.140 1.400 847.980 635.600 ;
    RECT 848.260 1.400 849.100 635.600 ;
    RECT 849.380 1.400 850.220 635.600 ;
    RECT 850.500 1.400 851.340 635.600 ;
    RECT 851.620 1.400 852.460 635.600 ;
    RECT 852.740 1.400 853.580 635.600 ;
    RECT 853.860 1.400 854.700 635.600 ;
    RECT 854.980 1.400 855.820 635.600 ;
    RECT 856.100 1.400 856.940 635.600 ;
    RECT 857.220 1.400 858.060 635.600 ;
    RECT 858.340 1.400 859.180 635.600 ;
    RECT 859.460 1.400 860.300 635.600 ;
    RECT 860.580 1.400 861.420 635.600 ;
    RECT 861.700 1.400 862.540 635.600 ;
    RECT 862.820 1.400 863.660 635.600 ;
    RECT 863.940 1.400 864.780 635.600 ;
    RECT 865.060 1.400 865.900 635.600 ;
    RECT 866.180 1.400 867.020 635.600 ;
    RECT 867.300 1.400 868.140 635.600 ;
    RECT 868.420 1.400 869.260 635.600 ;
    RECT 869.540 1.400 870.380 635.600 ;
    RECT 870.660 1.400 871.500 635.600 ;
    RECT 871.780 1.400 872.620 635.600 ;
    RECT 872.900 1.400 873.740 635.600 ;
    RECT 874.020 1.400 874.860 635.600 ;
    RECT 875.140 1.400 875.980 635.600 ;
    RECT 876.260 1.400 877.100 635.600 ;
    RECT 877.380 1.400 878.220 635.600 ;
    RECT 878.500 1.400 879.340 635.600 ;
    RECT 879.620 1.400 880.460 635.600 ;
    RECT 880.740 1.400 881.580 635.600 ;
    RECT 881.860 1.400 882.700 635.600 ;
    RECT 882.980 1.400 883.820 635.600 ;
    RECT 884.100 1.400 884.940 635.600 ;
    RECT 885.220 1.400 886.060 635.600 ;
    RECT 886.340 1.400 887.180 635.600 ;
    RECT 887.460 1.400 888.300 635.600 ;
    RECT 888.580 1.400 889.420 635.600 ;
    RECT 889.700 1.400 890.540 635.600 ;
    RECT 890.820 1.400 891.660 635.600 ;
    RECT 891.940 1.400 892.780 635.600 ;
    RECT 893.060 1.400 893.900 635.600 ;
    RECT 894.180 1.400 895.020 635.600 ;
    RECT 895.300 1.400 896.140 635.600 ;
    RECT 896.420 1.400 897.260 635.600 ;
    RECT 897.540 1.400 898.380 635.600 ;
    RECT 898.660 1.400 899.500 635.600 ;
    RECT 899.780 1.400 900.620 635.600 ;
    RECT 900.900 1.400 901.740 635.600 ;
    RECT 902.020 1.400 902.860 635.600 ;
    RECT 903.140 1.400 903.980 635.600 ;
    RECT 904.260 1.400 905.100 635.600 ;
    RECT 905.380 1.400 906.220 635.600 ;
    RECT 906.500 1.400 907.340 635.600 ;
    RECT 907.620 1.400 908.460 635.600 ;
    RECT 908.740 1.400 909.580 635.600 ;
    RECT 909.860 1.400 910.700 635.600 ;
    RECT 910.980 1.400 911.820 635.600 ;
    RECT 912.100 1.400 912.940 635.600 ;
    RECT 913.220 1.400 914.060 635.600 ;
    RECT 914.340 1.400 915.180 635.600 ;
    RECT 915.460 1.400 916.300 635.600 ;
    RECT 916.580 1.400 917.420 635.600 ;
    RECT 917.700 1.400 918.540 635.600 ;
    RECT 918.820 1.400 919.660 635.600 ;
    RECT 919.940 1.400 920.780 635.600 ;
    RECT 921.060 1.400 921.900 635.600 ;
    RECT 922.180 1.400 923.020 635.600 ;
    RECT 923.300 1.400 924.140 635.600 ;
    RECT 924.420 1.400 925.260 635.600 ;
    RECT 925.540 1.400 926.380 635.600 ;
    RECT 926.660 1.400 927.500 635.600 ;
    RECT 927.780 1.400 928.620 635.600 ;
    RECT 928.900 1.400 929.740 635.600 ;
    RECT 930.020 1.400 930.860 635.600 ;
    RECT 931.140 1.400 931.980 635.600 ;
    RECT 932.260 1.400 933.100 635.600 ;
    RECT 933.380 1.400 934.220 635.600 ;
    RECT 934.500 1.400 935.340 635.600 ;
    RECT 935.620 1.400 936.460 635.600 ;
    RECT 936.740 1.400 937.580 635.600 ;
    RECT 937.860 1.400 938.700 635.600 ;
    RECT 938.980 1.400 939.820 635.600 ;
    RECT 940.100 1.400 940.940 635.600 ;
    RECT 941.220 1.400 942.060 635.600 ;
    RECT 942.340 1.400 943.180 635.600 ;
    RECT 943.460 1.400 944.300 635.600 ;
    RECT 944.580 1.400 945.420 635.600 ;
    RECT 945.700 1.400 946.540 635.600 ;
    RECT 946.820 1.400 947.660 635.600 ;
    RECT 947.940 1.400 948.780 635.600 ;
    RECT 949.060 1.400 949.900 635.600 ;
    RECT 950.180 1.400 951.020 635.600 ;
    RECT 951.300 1.400 952.140 635.600 ;
    RECT 952.420 1.400 953.260 635.600 ;
    RECT 953.540 1.400 954.380 635.600 ;
    RECT 954.660 1.400 955.500 635.600 ;
    RECT 955.780 1.400 956.620 635.600 ;
    RECT 956.900 1.400 957.740 635.600 ;
    RECT 958.020 1.400 958.860 635.600 ;
    RECT 959.140 1.400 959.980 635.600 ;
    RECT 960.260 1.400 961.100 635.600 ;
    RECT 961.380 1.400 962.220 635.600 ;
    RECT 962.500 1.400 963.340 635.600 ;
    RECT 963.620 1.400 964.460 635.600 ;
    RECT 964.740 1.400 965.580 635.600 ;
    RECT 965.860 1.400 966.700 635.600 ;
    RECT 966.980 1.400 967.820 635.600 ;
    RECT 968.100 1.400 968.940 635.600 ;
    RECT 969.220 1.400 970.060 635.600 ;
    RECT 970.340 1.400 971.180 635.600 ;
    RECT 971.460 1.400 972.300 635.600 ;
    RECT 972.580 1.400 973.420 635.600 ;
    RECT 973.700 1.400 974.540 635.600 ;
    RECT 974.820 1.400 975.660 635.600 ;
    RECT 975.940 1.400 976.780 635.600 ;
    RECT 977.060 1.400 977.900 635.600 ;
    RECT 978.180 1.400 979.020 635.600 ;
    RECT 979.300 1.400 980.140 635.600 ;
    RECT 980.420 1.400 981.260 635.600 ;
    RECT 981.540 1.400 982.380 635.600 ;
    RECT 982.660 1.400 983.500 635.600 ;
    RECT 983.780 1.400 984.620 635.600 ;
    RECT 984.900 1.400 985.740 635.600 ;
    RECT 986.020 1.400 986.860 635.600 ;
    RECT 987.140 1.400 987.980 635.600 ;
    RECT 988.260 1.400 989.100 635.600 ;
    RECT 989.380 1.400 990.220 635.600 ;
    RECT 990.500 1.400 991.340 635.600 ;
    RECT 991.620 1.400 992.460 635.600 ;
    RECT 992.740 1.400 993.580 635.600 ;
    RECT 993.860 1.400 994.700 635.600 ;
    RECT 994.980 1.400 995.820 635.600 ;
    RECT 996.100 1.400 996.940 635.600 ;
    RECT 997.220 1.400 998.060 635.600 ;
    RECT 998.340 1.400 999.180 635.600 ;
    RECT 999.460 1.400 1000.300 635.600 ;
    RECT 1000.580 1.400 1001.420 635.600 ;
    RECT 1001.700 1.400 1002.540 635.600 ;
    RECT 1002.820 1.400 1003.660 635.600 ;
    RECT 1003.940 1.400 1004.780 635.600 ;
    RECT 1005.060 1.400 1005.900 635.600 ;
    RECT 1006.180 1.400 1007.020 635.600 ;
    RECT 1007.300 1.400 1008.140 635.600 ;
    RECT 1008.420 1.400 1009.260 635.600 ;
    RECT 1009.540 1.400 1010.380 635.600 ;
    RECT 1010.660 1.400 1011.500 635.600 ;
    RECT 1011.780 1.400 1012.620 635.600 ;
    RECT 1012.900 1.400 1013.740 635.600 ;
    RECT 1014.020 1.400 1014.860 635.600 ;
    RECT 1015.140 1.400 1015.980 635.600 ;
    RECT 1016.260 1.400 1017.100 635.600 ;
    RECT 1017.380 1.400 1018.220 635.600 ;
    RECT 1018.500 1.400 1019.340 635.600 ;
    RECT 1019.620 1.400 1020.460 635.600 ;
    RECT 1020.740 1.400 1021.580 635.600 ;
    RECT 1021.860 1.400 1022.700 635.600 ;
    RECT 1022.980 1.400 1023.820 635.600 ;
    RECT 1024.100 1.400 1024.940 635.600 ;
    RECT 1025.220 1.400 1026.060 635.600 ;
    RECT 1026.340 1.400 1027.180 635.600 ;
    RECT 1027.460 1.400 1028.300 635.600 ;
    RECT 1028.580 1.400 1029.420 635.600 ;
    RECT 1029.700 1.400 1030.540 635.600 ;
    RECT 1030.820 1.400 1031.660 635.600 ;
    RECT 1031.940 1.400 1032.780 635.600 ;
    RECT 1033.060 1.400 1033.900 635.600 ;
    RECT 1034.180 1.400 1035.020 635.600 ;
    RECT 1035.300 1.400 1036.140 635.600 ;
    RECT 1036.420 1.400 1037.260 635.600 ;
    RECT 1037.540 1.400 1038.380 635.600 ;
    RECT 1038.660 1.400 1039.500 635.600 ;
    RECT 1039.780 1.400 1040.620 635.600 ;
    RECT 1040.900 1.400 1041.740 635.600 ;
    RECT 1042.020 1.400 1042.860 635.600 ;
    RECT 1043.140 1.400 1043.980 635.600 ;
    RECT 1044.260 1.400 1045.100 635.600 ;
    RECT 1045.380 1.400 1046.220 635.600 ;
    RECT 1046.500 1.400 1047.340 635.600 ;
    RECT 1047.620 1.400 1048.460 635.600 ;
    RECT 1048.740 1.400 1049.580 635.600 ;
    RECT 1049.860 1.400 1050.700 635.600 ;
    RECT 1050.980 1.400 1051.820 635.600 ;
    RECT 1052.100 1.400 1052.940 635.600 ;
    RECT 1053.220 1.400 1054.060 635.600 ;
    RECT 1054.340 1.400 1055.180 635.600 ;
    RECT 1055.460 1.400 1056.300 635.600 ;
    RECT 1056.580 1.400 1057.420 635.600 ;
    RECT 1057.700 1.400 1058.540 635.600 ;
    RECT 1058.820 1.400 1059.660 635.600 ;
    RECT 1059.940 1.400 1060.780 635.600 ;
    RECT 1061.060 1.400 1061.900 635.600 ;
    RECT 1062.180 1.400 1063.020 635.600 ;
    RECT 1063.300 1.400 1064.140 635.600 ;
    RECT 1064.420 1.400 1065.260 635.600 ;
    RECT 1065.540 1.400 1066.380 635.600 ;
    RECT 1066.660 1.400 1067.500 635.600 ;
    RECT 1067.780 1.400 1068.620 635.600 ;
    RECT 1068.900 1.400 1069.740 635.600 ;
    RECT 1070.020 1.400 1070.860 635.600 ;
    RECT 1071.140 1.400 1071.980 635.600 ;
    RECT 1072.260 1.400 1073.100 635.600 ;
    RECT 1073.380 1.400 1074.220 635.600 ;
    RECT 1074.500 1.400 1075.340 635.600 ;
    RECT 1075.620 1.400 1076.460 635.600 ;
    RECT 1076.740 1.400 1077.580 635.600 ;
    RECT 1077.860 1.400 1078.700 635.600 ;
    RECT 1078.980 1.400 1079.820 635.600 ;
    RECT 1080.100 1.400 1080.940 635.600 ;
    RECT 1081.220 1.400 1082.060 635.600 ;
    RECT 1082.340 1.400 1083.180 635.600 ;
    RECT 1083.460 1.400 1084.300 635.600 ;
    RECT 1084.580 1.400 1085.420 635.600 ;
    RECT 1085.700 1.400 1086.540 635.600 ;
    RECT 1086.820 1.400 1087.660 635.600 ;
    RECT 1087.940 1.400 1088.780 635.600 ;
    RECT 1089.060 1.400 1089.900 635.600 ;
    RECT 1090.180 1.400 1091.020 635.600 ;
    RECT 1091.300 1.400 1092.140 635.600 ;
    RECT 1092.420 1.400 1093.260 635.600 ;
    RECT 1093.540 1.400 1094.380 635.600 ;
    RECT 1094.660 1.400 1095.500 635.600 ;
    RECT 1095.780 1.400 1096.620 635.600 ;
    RECT 1096.900 1.400 1097.740 635.600 ;
    RECT 1098.020 1.400 1098.860 635.600 ;
    RECT 1099.140 1.400 1099.980 635.600 ;
    RECT 1100.260 1.400 1101.100 635.600 ;
    RECT 1101.380 1.400 1102.220 635.600 ;
    RECT 1102.500 1.400 1103.340 635.600 ;
    RECT 1103.620 1.400 1104.460 635.600 ;
    RECT 1104.740 1.400 1105.580 635.600 ;
    RECT 1105.860 1.400 1106.700 635.600 ;
    RECT 1106.980 1.400 1107.820 635.600 ;
    RECT 1108.100 1.400 1108.940 635.600 ;
    RECT 1109.220 1.400 1110.060 635.600 ;
    RECT 1110.340 1.400 1111.180 635.600 ;
    RECT 1111.460 1.400 1112.300 635.600 ;
    RECT 1112.580 1.400 1113.420 635.600 ;
    RECT 1113.700 1.400 1114.540 635.600 ;
    RECT 1114.820 1.400 1115.660 635.600 ;
    RECT 1115.940 1.400 1116.780 635.600 ;
    RECT 1117.060 1.400 1117.900 635.600 ;
    RECT 1118.180 1.400 1119.020 635.600 ;
    RECT 1119.300 1.400 1120.140 635.600 ;
    RECT 1120.420 1.400 1121.260 635.600 ;
    RECT 1121.540 1.400 1122.380 635.600 ;
    RECT 1122.660 1.400 1123.500 635.600 ;
    RECT 1123.780 1.400 1124.620 635.600 ;
    RECT 1124.900 1.400 1125.740 635.600 ;
    RECT 1126.020 1.400 1126.860 635.600 ;
    RECT 1127.140 1.400 1127.980 635.600 ;
    RECT 1128.260 1.400 1129.100 635.600 ;
    RECT 1129.380 1.400 1130.220 635.600 ;
    RECT 1130.500 1.400 1131.340 635.600 ;
    RECT 1131.620 1.400 1132.460 635.600 ;
    RECT 1132.740 1.400 1133.580 635.600 ;
    RECT 1133.860 1.400 1134.700 635.600 ;
    RECT 1134.980 1.400 1135.820 635.600 ;
    RECT 1136.100 1.400 1136.940 635.600 ;
    RECT 1137.220 1.400 1138.060 635.600 ;
    RECT 1138.340 1.400 1139.180 635.600 ;
    RECT 1139.460 1.400 1140.300 635.600 ;
    RECT 1140.580 1.400 1141.420 635.600 ;
    RECT 1141.700 1.400 1142.540 635.600 ;
    RECT 1142.820 1.400 1143.660 635.600 ;
    RECT 1143.940 1.400 1144.780 635.600 ;
    RECT 1145.060 1.400 1145.900 635.600 ;
    RECT 1146.180 1.400 1147.020 635.600 ;
    RECT 1147.300 1.400 1148.140 635.600 ;
    RECT 1148.420 1.400 1149.260 635.600 ;
    RECT 1149.540 1.400 1150.380 635.600 ;
    RECT 1150.660 1.400 1151.500 635.600 ;
    RECT 1151.780 1.400 1152.620 635.600 ;
    RECT 1152.900 1.400 1153.740 635.600 ;
    RECT 1154.020 1.400 1154.860 635.600 ;
    RECT 1155.140 1.400 1155.980 635.600 ;
    RECT 1156.260 1.400 1157.100 635.600 ;
    RECT 1157.380 1.400 1158.220 635.600 ;
    RECT 1158.500 1.400 1159.340 635.600 ;
    RECT 1159.620 1.400 1160.460 635.600 ;
    RECT 1160.740 1.400 1161.580 635.600 ;
    RECT 1161.860 1.400 1162.700 635.600 ;
    RECT 1162.980 1.400 1163.820 635.600 ;
    RECT 1164.100 1.400 1164.940 635.600 ;
    RECT 1165.220 1.400 1166.060 635.600 ;
    RECT 1166.340 1.400 1167.180 635.600 ;
    RECT 1167.460 1.400 1168.300 635.600 ;
    RECT 1168.580 1.400 1169.420 635.600 ;
    RECT 1169.700 1.400 1170.540 635.600 ;
    RECT 1170.820 1.400 1171.660 635.600 ;
    RECT 1171.940 1.400 1172.780 635.600 ;
    RECT 1173.060 1.400 1173.900 635.600 ;
    RECT 1174.180 1.400 1175.020 635.600 ;
    RECT 1175.300 1.400 1176.140 635.600 ;
    RECT 1176.420 1.400 1177.260 635.600 ;
    RECT 1177.540 1.400 1178.380 635.600 ;
    RECT 1178.660 1.400 1179.500 635.600 ;
    RECT 1179.780 1.400 1180.620 635.600 ;
    RECT 1180.900 1.400 1181.740 635.600 ;
    RECT 1182.020 1.400 1182.860 635.600 ;
    RECT 1183.140 1.400 1183.980 635.600 ;
    RECT 1184.260 1.400 1185.100 635.600 ;
    RECT 1185.380 1.400 1186.220 635.600 ;
    RECT 1186.500 1.400 1187.340 635.600 ;
    RECT 1187.620 1.400 1188.460 635.600 ;
    RECT 1188.740 1.400 1189.580 635.600 ;
    RECT 1189.860 1.400 1190.700 635.600 ;
    RECT 1190.980 1.400 1191.820 635.600 ;
    RECT 1192.100 1.400 1192.940 635.600 ;
    RECT 1193.220 1.400 1194.060 635.600 ;
    RECT 1194.340 1.400 1195.180 635.600 ;
    RECT 1195.460 1.400 1196.300 635.600 ;
    RECT 1196.580 1.400 1197.420 635.600 ;
    RECT 1197.700 1.400 1198.540 635.600 ;
    RECT 1198.820 1.400 1199.660 635.600 ;
    RECT 1199.940 1.400 1200.780 635.600 ;
    RECT 1201.060 1.400 1201.900 635.600 ;
    RECT 1202.180 1.400 1203.020 635.600 ;
    RECT 1203.300 1.400 1204.140 635.600 ;
    RECT 1204.420 1.400 1205.260 635.600 ;
    RECT 1205.540 1.400 1206.380 635.600 ;
    RECT 1206.660 1.400 1207.500 635.600 ;
    RECT 1207.780 1.400 1208.620 635.600 ;
    RECT 1208.900 1.400 1209.740 635.600 ;
    RECT 1210.020 1.400 1210.860 635.600 ;
    RECT 1211.140 1.400 1211.980 635.600 ;
    RECT 1212.260 1.400 1213.100 635.600 ;
    RECT 1213.380 1.400 1214.220 635.600 ;
    RECT 1214.500 1.400 1215.340 635.600 ;
    RECT 1215.620 1.400 1216.460 635.600 ;
    RECT 1216.740 1.400 1217.580 635.600 ;
    RECT 1217.860 1.400 1218.700 635.600 ;
    RECT 1218.980 1.400 1219.820 635.600 ;
    RECT 1220.100 1.400 1220.940 635.600 ;
    RECT 1221.220 1.400 1222.060 635.600 ;
    RECT 1222.340 1.400 1223.180 635.600 ;
    RECT 1223.460 1.400 1224.300 635.600 ;
    RECT 1224.580 1.400 1225.420 635.600 ;
    RECT 1225.700 1.400 1226.540 635.600 ;
    RECT 1226.820 1.400 1227.660 635.600 ;
    RECT 1227.940 1.400 1228.780 635.600 ;
    RECT 1229.060 1.400 1229.900 635.600 ;
    RECT 1230.180 1.400 1231.020 635.600 ;
    RECT 1231.300 1.400 1232.140 635.600 ;
    RECT 1232.420 1.400 1233.260 635.600 ;
    RECT 1233.540 1.400 1234.380 635.600 ;
    RECT 1234.660 1.400 1235.500 635.600 ;
    RECT 1235.780 1.400 1236.620 635.600 ;
    RECT 1236.900 1.400 1237.740 635.600 ;
    RECT 1238.020 1.400 1238.860 635.600 ;
    RECT 1239.140 1.400 1239.980 635.600 ;
    RECT 1240.260 1.400 1241.100 635.600 ;
    RECT 1241.380 1.400 1242.220 635.600 ;
    RECT 1242.500 1.400 1243.340 635.600 ;
    RECT 1243.620 1.400 1244.460 635.600 ;
    RECT 1244.740 1.400 1245.580 635.600 ;
    RECT 1245.860 1.400 1246.700 635.600 ;
    RECT 1246.980 1.400 1247.820 635.600 ;
    RECT 1248.100 1.400 1248.940 635.600 ;
    RECT 1249.220 1.400 1250.060 635.600 ;
    RECT 1250.340 1.400 1251.180 635.600 ;
    RECT 1251.460 1.400 1252.300 635.600 ;
    RECT 1252.580 1.400 1253.420 635.600 ;
    RECT 1253.700 1.400 1254.540 635.600 ;
    RECT 1254.820 1.400 1255.660 635.600 ;
    RECT 1255.940 1.400 1256.780 635.600 ;
    RECT 1257.060 1.400 1257.900 635.600 ;
    RECT 1258.180 1.400 1259.020 635.600 ;
    RECT 1259.300 1.400 1260.140 635.600 ;
    RECT 1260.420 1.400 1261.260 635.600 ;
    RECT 1261.540 1.400 1262.380 635.600 ;
    RECT 1262.660 1.400 1263.500 635.600 ;
    RECT 1263.780 1.400 1264.620 635.600 ;
    RECT 1264.900 1.400 1265.740 635.600 ;
    RECT 1266.020 1.400 1266.860 635.600 ;
    RECT 1267.140 1.400 1267.980 635.600 ;
    RECT 1268.260 1.400 1269.100 635.600 ;
    RECT 1269.380 1.400 1270.220 635.600 ;
    RECT 1270.500 1.400 1271.340 635.600 ;
    RECT 1271.620 1.400 1272.460 635.600 ;
    RECT 1272.740 1.400 1273.580 635.600 ;
    RECT 1273.860 1.400 1274.700 635.600 ;
    RECT 1274.980 1.400 1275.820 635.600 ;
    RECT 1276.100 1.400 1276.940 635.600 ;
    RECT 1277.220 1.400 1278.060 635.600 ;
    RECT 1278.340 1.400 1279.180 635.600 ;
    RECT 1279.460 1.400 1280.300 635.600 ;
    RECT 1280.580 1.400 1281.420 635.600 ;
    RECT 1281.700 1.400 1282.540 635.600 ;
    RECT 1282.820 1.400 1283.660 635.600 ;
    RECT 1283.940 1.400 1284.780 635.600 ;
    RECT 1285.060 1.400 1285.900 635.600 ;
    RECT 1286.180 1.400 1287.020 635.600 ;
    RECT 1287.300 1.400 1288.140 635.600 ;
    RECT 1288.420 1.400 1289.260 635.600 ;
    RECT 1289.540 1.400 1290.380 635.600 ;
    RECT 1290.660 1.400 1291.500 635.600 ;
    RECT 1291.780 1.400 1292.620 635.600 ;
    RECT 1292.900 1.400 1293.740 635.600 ;
    RECT 1294.020 1.400 1294.860 635.600 ;
    RECT 1295.140 1.400 1295.980 635.600 ;
    RECT 1296.260 1.400 1297.100 635.600 ;
    RECT 1297.380 1.400 1298.220 635.600 ;
    RECT 1298.500 1.400 1299.340 635.600 ;
    RECT 1299.620 1.400 1300.460 635.600 ;
    RECT 1300.740 1.400 1301.580 635.600 ;
    RECT 1301.860 1.400 1302.700 635.600 ;
    RECT 1302.980 1.400 1303.820 635.600 ;
    RECT 1304.100 1.400 1304.940 635.600 ;
    RECT 1305.220 1.400 1306.060 635.600 ;
    RECT 1306.340 1.400 1307.180 635.600 ;
    RECT 1307.460 1.400 1308.300 635.600 ;
    RECT 1308.580 1.400 1309.420 635.600 ;
    RECT 1309.700 1.400 1310.540 635.600 ;
    RECT 1310.820 1.400 1311.660 635.600 ;
    RECT 1311.940 1.400 1312.780 635.600 ;
    RECT 1313.060 1.400 1313.900 635.600 ;
    RECT 1314.180 1.400 1315.020 635.600 ;
    RECT 1315.300 1.400 1316.140 635.600 ;
    RECT 1316.420 1.400 1317.260 635.600 ;
    RECT 1317.540 1.400 1318.380 635.600 ;
    RECT 1318.660 1.400 1319.500 635.600 ;
    RECT 1319.780 1.400 1320.620 635.600 ;
    RECT 1320.900 1.400 1321.740 635.600 ;
    RECT 1322.020 1.400 1322.860 635.600 ;
    RECT 1323.140 1.400 1323.980 635.600 ;
    RECT 1324.260 1.400 1325.100 635.600 ;
    RECT 1325.380 1.400 1326.220 635.600 ;
    RECT 1326.500 1.400 1327.340 635.600 ;
    RECT 1327.620 1.400 1328.460 635.600 ;
    RECT 1328.740 1.400 1329.580 635.600 ;
    RECT 1329.860 1.400 1330.700 635.600 ;
    RECT 1330.980 1.400 1331.820 635.600 ;
    RECT 1332.100 1.400 1332.940 635.600 ;
    RECT 1333.220 1.400 1334.060 635.600 ;
    RECT 1334.340 1.400 1335.180 635.600 ;
    RECT 1335.460 1.400 1336.300 635.600 ;
    RECT 1336.580 1.400 1337.420 635.600 ;
    RECT 1337.700 1.400 1338.540 635.600 ;
    RECT 1338.820 1.400 1339.660 635.600 ;
    RECT 1339.940 1.400 1340.780 635.600 ;
    RECT 1341.060 1.400 1341.900 635.600 ;
    RECT 1342.180 1.400 1343.020 635.600 ;
    RECT 1343.300 1.400 1344.140 635.600 ;
    RECT 1344.420 1.400 1345.260 635.600 ;
    RECT 1345.540 1.400 1346.380 635.600 ;
    RECT 1346.660 1.400 1347.500 635.600 ;
    RECT 1347.780 1.400 1348.620 635.600 ;
    RECT 1348.900 1.400 1349.740 635.600 ;
    RECT 1350.020 1.400 1350.860 635.600 ;
    RECT 1351.140 1.400 1351.980 635.600 ;
    RECT 1352.260 1.400 1353.100 635.600 ;
    RECT 1353.380 1.400 1354.220 635.600 ;
    RECT 1354.500 1.400 1355.340 635.600 ;
    RECT 1355.620 1.400 1356.460 635.600 ;
    RECT 1356.740 1.400 1357.580 635.600 ;
    RECT 1357.860 1.400 1358.700 635.600 ;
    RECT 1358.980 1.400 1359.820 635.600 ;
    RECT 1360.100 1.400 1360.940 635.600 ;
    RECT 1361.220 1.400 1362.060 635.600 ;
    RECT 1362.340 1.400 1363.180 635.600 ;
    RECT 1363.460 1.400 1364.300 635.600 ;
    RECT 1364.580 1.400 1365.420 635.600 ;
    RECT 1365.700 1.400 1366.540 635.600 ;
    RECT 1366.820 1.400 1367.660 635.600 ;
    RECT 1367.940 1.400 1368.780 635.600 ;
    RECT 1369.060 1.400 1369.900 635.600 ;
    RECT 1370.180 1.400 1371.020 635.600 ;
    RECT 1371.300 1.400 1372.140 635.600 ;
    RECT 1372.420 1.400 1373.260 635.600 ;
    RECT 1373.540 1.400 1374.380 635.600 ;
    RECT 1374.660 1.400 1375.500 635.600 ;
    RECT 1375.780 1.400 1376.620 635.600 ;
    RECT 1376.900 1.400 1377.740 635.600 ;
    RECT 1378.020 1.400 1378.860 635.600 ;
    RECT 1379.140 1.400 1379.980 635.600 ;
    RECT 1380.260 1.400 1381.100 635.600 ;
    RECT 1381.380 1.400 1382.220 635.600 ;
    RECT 1382.500 1.400 1383.340 635.600 ;
    RECT 1383.620 1.400 1384.460 635.600 ;
    RECT 1384.740 1.400 1385.580 635.600 ;
    RECT 1385.860 1.400 1386.700 635.600 ;
    RECT 1386.980 1.400 1387.820 635.600 ;
    RECT 1388.100 1.400 1388.940 635.600 ;
    RECT 1389.220 1.400 1390.060 635.600 ;
    RECT 1390.340 1.400 1391.180 635.600 ;
    RECT 1391.460 1.400 1392.300 635.600 ;
    RECT 1392.580 1.400 1393.420 635.600 ;
    RECT 1393.700 1.400 1394.540 635.600 ;
    RECT 1394.820 1.400 1395.660 635.600 ;
    RECT 1395.940 1.400 1396.780 635.600 ;
    RECT 1397.060 1.400 1397.900 635.600 ;
    RECT 1398.180 1.400 1399.020 635.600 ;
    RECT 1399.300 1.400 1400.140 635.600 ;
    RECT 1400.420 1.400 1401.260 635.600 ;
    RECT 1401.540 1.400 1402.380 635.600 ;
    RECT 1402.660 1.400 1403.500 635.600 ;
    RECT 1403.780 1.400 1404.620 635.600 ;
    RECT 1404.900 1.400 1405.740 635.600 ;
    RECT 1406.020 1.400 1406.860 635.600 ;
    RECT 1407.140 1.400 1407.980 635.600 ;
    RECT 1408.260 1.400 1409.100 635.600 ;
    RECT 1409.380 1.400 1410.220 635.600 ;
    RECT 1410.500 1.400 1411.340 635.600 ;
    RECT 1411.620 1.400 1412.460 635.600 ;
    RECT 1412.740 1.400 1413.580 635.600 ;
    RECT 1413.860 1.400 1414.700 635.600 ;
    RECT 1414.980 1.400 1415.820 635.600 ;
    RECT 1416.100 1.400 1416.940 635.600 ;
    RECT 1417.220 1.400 1418.060 635.600 ;
    RECT 1418.340 1.400 1419.180 635.600 ;
    RECT 1419.460 1.400 1420.300 635.600 ;
    RECT 1420.580 1.400 1421.420 635.600 ;
    RECT 1421.700 1.400 1422.540 635.600 ;
    RECT 1422.820 1.400 1423.660 635.600 ;
    RECT 1423.940 1.400 1424.780 635.600 ;
    RECT 1425.060 1.400 1425.900 635.600 ;
    RECT 1426.180 1.400 1427.020 635.600 ;
    RECT 1427.300 1.400 1428.140 635.600 ;
    RECT 1428.420 1.400 1429.260 635.600 ;
    RECT 1429.540 1.400 1430.380 635.600 ;
    RECT 1430.660 1.400 1431.500 635.600 ;
    RECT 1431.780 1.400 1432.620 635.600 ;
    RECT 1432.900 1.400 1433.740 635.600 ;
    RECT 1434.020 1.400 1434.860 635.600 ;
    RECT 1435.140 1.400 1435.980 635.600 ;
    RECT 1436.260 1.400 1437.100 635.600 ;
    RECT 1437.380 1.400 1438.220 635.600 ;
    RECT 1438.500 1.400 1439.340 635.600 ;
    RECT 1439.620 1.400 1440.460 635.600 ;
    RECT 1440.740 1.400 1441.580 635.600 ;
    RECT 1441.860 1.400 1442.700 635.600 ;
    RECT 1442.980 1.400 1443.820 635.600 ;
    RECT 1444.100 1.400 1444.940 635.600 ;
    RECT 1445.220 1.400 1446.060 635.600 ;
    RECT 1446.340 1.400 1447.180 635.600 ;
    RECT 1447.460 1.400 1448.300 635.600 ;
    RECT 1448.580 1.400 1449.420 635.600 ;
    RECT 1449.700 1.400 1450.540 635.600 ;
    RECT 1450.820 1.400 1451.660 635.600 ;
    RECT 1451.940 1.400 1452.780 635.600 ;
    RECT 1453.060 1.400 1453.900 635.600 ;
    RECT 1454.180 1.400 1455.020 635.600 ;
    RECT 1455.300 1.400 1456.140 635.600 ;
    RECT 1456.420 1.400 1457.260 635.600 ;
    RECT 1457.540 1.400 1458.380 635.600 ;
    RECT 1458.660 1.400 1459.500 635.600 ;
    RECT 1459.780 1.400 1461.480 635.600 ;
    LAYER OVERLAP ;
    RECT 0 0 1461.480 637.000 ;
  END
END sram_64x16384_1rw

END LIBRARY
